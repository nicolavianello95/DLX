
module SNPS_CLOCK_GATE_HIGH_HDU ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19519, net19521, net19523, net19524, net19527, net19530;
  assign net19519 = EN;
  assign net19521 = CLK;
  assign ENCLK = net19523;
  assign net19530 = TE;

  DLL_X1 latch ( .D(net19524), .GN(net19521), .Q(net19527) );
  AND2_X1 main_gate ( .A1(net19527), .A2(net19521), .ZN(net19523) );
  OR2_X1 test_or ( .A1(net19519), .A2(net19530), .ZN(net19524) );
endmodule


module HDU ( INSTR_ID, INSTR_EXE, .HDU_OUTS({\HDU_OUTS[PC_EN] , 
        \HDU_OUTS[IF_EN] , \HDU_OUTS[ID_EN] , \HDU_OUTS[EXE_EN] , 
        \HDU_OUTS[MEM_EN] , \HDU_OUTS[WB_EN] , \HDU_OUTS[ID_BUBBLE] , 
        \HDU_OUTS[EXE_BUBBLE] , \HDU_OUTS[MEM_BUBBLE] , \HDU_OUTS[WB_BUBBLE] }
        ), clk, rst, misprediction_BAR );
  input [31:0] INSTR_ID;
  input [31:0] INSTR_EXE;
  input clk, rst, misprediction_BAR;
  output \HDU_OUTS[PC_EN] , \HDU_OUTS[IF_EN] , \HDU_OUTS[ID_EN] ,
         \HDU_OUTS[EXE_EN] , \HDU_OUTS[MEM_EN] , \HDU_OUTS[WB_EN] ,
         \HDU_OUTS[ID_BUBBLE] , \HDU_OUTS[EXE_BUBBLE] , \HDU_OUTS[MEM_BUBBLE] ,
         \HDU_OUTS[WB_BUBBLE] ;
  wire   INSTR_EXE_31, INSTR_EXE_30, INSTR_EXE_29, INSTR_EXE_28, INSTR_EXE_27,
         INSTR_EXE_26, INSTR_EXE_5, INSTR_EXE_4, INSTR_EXE_3, INSTR_EXE_2,
         INSTR_EXE_1, INSTR_EXE_0, misprediction, \HDU_OUTS[PC_EN] , N683,
         N689, net19535, n5, n6, n1, n2, n3, n4, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39;
  assign INSTR_EXE_31 = INSTR_EXE[31];
  assign INSTR_EXE_30 = INSTR_EXE[30];
  assign INSTR_EXE_29 = INSTR_EXE[29];
  assign INSTR_EXE_28 = INSTR_EXE[28];
  assign INSTR_EXE_27 = INSTR_EXE[27];
  assign INSTR_EXE_26 = INSTR_EXE[26];
  assign INSTR_EXE_5 = INSTR_EXE[5];
  assign INSTR_EXE_4 = INSTR_EXE[4];
  assign INSTR_EXE_3 = INSTR_EXE[3];
  assign INSTR_EXE_2 = INSTR_EXE[2];
  assign INSTR_EXE_1 = INSTR_EXE[1];
  assign INSTR_EXE_0 = INSTR_EXE[0];
  assign misprediction = misprediction_BAR;
  assign \HDU_OUTS[ID_EN]  = \HDU_OUTS[PC_EN] ;

  SNPS_CLOCK_GATE_HIGH_HDU clk_gate_count_reg ( .CLK(clk), .EN(N683), .ENCLK(
        net19535), .TE(1'b0) );
  DFFR_X1 \count_reg[0]  ( .D(n6), .CK(net19535), .RN(rst), .QN(n6) );
  DFFR_X1 \count_reg[1]  ( .D(N689), .CK(net19535), .RN(rst), .QN(n5) );
  OR2_X1 U3 ( .A1(n1), .A2(n37), .ZN(n2) );
  NAND4_X1 U4 ( .A1(n25), .A2(n26), .A3(n27), .A4(n28), .ZN(n3) );
  NOR3_X1 U5 ( .A1(INSTR_ID[28]), .A2(INSTR_ID[29]), .A3(INSTR_ID[31]), .ZN(n4) );
  NAND2_X1 U6 ( .A1(INSTR_ID[27]), .A2(n4), .ZN(n7) );
  OAI22_X1 U7 ( .A1(INSTR_EXE[17]), .A2(n3), .B1(INSTR_ID[30]), .B2(n7), .ZN(
        n8) );
  INV_X1 U8 ( .A(INSTR_EXE_26), .ZN(n1) );
  AOI221_X1 U9 ( .B1(INSTR_EXE_28), .B2(INSTR_EXE_27), .C1(n1), .C2(
        INSTR_EXE_27), .A(INSTR_EXE_30), .ZN(n9) );
  INV_X1 U10 ( .A(INSTR_EXE[17]), .ZN(n10) );
  OAI22_X1 U11 ( .A1(n10), .A2(INSTR_ID[22]), .B1(n25), .B2(INSTR_ID[25]), 
        .ZN(n11) );
  AOI221_X1 U12 ( .B1(n10), .B2(INSTR_ID[22]), .C1(INSTR_ID[25]), .C2(n25), 
        .A(n11), .ZN(n12) );
  OAI22_X1 U13 ( .A1(n26), .A2(INSTR_ID[21]), .B1(n27), .B2(INSTR_ID[24]), 
        .ZN(n13) );
  AOI221_X1 U14 ( .B1(n26), .B2(INSTR_ID[21]), .C1(INSTR_ID[24]), .C2(n27), 
        .A(n13), .ZN(n14) );
  OAI211_X1 U15 ( .C1(n28), .C2(INSTR_ID[23]), .A(n14), .B(n12), .ZN(n15) );
  AOI21_X1 U16 ( .B1(n28), .B2(INSTR_ID[23]), .A(n15), .ZN(n16) );
  AOI22_X1 U17 ( .A1(n27), .A2(INSTR_ID[19]), .B1(n26), .B2(INSTR_ID[16]), 
        .ZN(n17) );
  OAI221_X1 U18 ( .B1(n27), .B2(INSTR_ID[19]), .C1(n26), .C2(INSTR_ID[16]), 
        .A(n17), .ZN(n18) );
  AOI21_X1 U19 ( .B1(n25), .B2(INSTR_ID[20]), .A(INSTR_ID[26]), .ZN(n19) );
  OAI211_X1 U20 ( .C1(n25), .C2(INSTR_ID[20]), .A(n4), .B(n19), .ZN(n20) );
  AOI22_X1 U21 ( .A1(n28), .A2(INSTR_ID[18]), .B1(n10), .B2(INSTR_ID[17]), 
        .ZN(n21) );
  OAI221_X1 U22 ( .B1(n28), .B2(INSTR_ID[18]), .C1(n10), .C2(INSTR_ID[17]), 
        .A(n21), .ZN(n22) );
  NOR4_X1 U23 ( .A1(INSTR_ID[30]), .A2(n18), .A3(n20), .A4(n22), .ZN(n23) );
  OAI22_X1 U24 ( .A1(n36), .A2(n9), .B1(n16), .B2(n23), .ZN(n24) );
  AOI211_X1 U25 ( .C1(n36), .C2(n2), .A(n8), .B(n24), .ZN(
        \HDU_OUTS[EXE_BUBBLE] ) );
  XOR2_X1 U26 ( .A(n6), .B(n5), .Z(N689) );
  NOR2_X1 U27 ( .A1(\HDU_OUTS[EXE_BUBBLE] ), .A2(\HDU_OUTS[MEM_BUBBLE] ), .ZN(
        \HDU_OUTS[PC_EN] ) );
  INV_X1 U28 ( .A(\HDU_OUTS[EXE_EN] ), .ZN(\HDU_OUTS[MEM_BUBBLE] ) );
  OAI21_X1 U29 ( .B1(n5), .B2(n6), .A(N683), .ZN(\HDU_OUTS[EXE_EN] ) );
  OR4_X1 U30 ( .A1(INSTR_EXE_0), .A2(INSTR_EXE_5), .A3(n34), .A4(n33), .ZN(n35) );
  AND2_X1 U31 ( .A1(\HDU_OUTS[PC_EN] ), .A2(misprediction), .ZN(
        \HDU_OUTS[IF_EN] ) );
  NOR2_X1 U32 ( .A1(misprediction), .A2(n39), .ZN(\HDU_OUTS[ID_BUBBLE] ) );
  OR4_X1 U33 ( .A1(INSTR_EXE_30), .A2(INSTR_EXE_29), .A3(INSTR_EXE_27), .A4(
        INSTR_EXE_28), .ZN(n34) );
  INV_X1 U34 ( .A(INSTR_EXE_29), .ZN(n29) );
  OAI21_X1 U35 ( .B1(INSTR_EXE_30), .B2(n29), .A(INSTR_EXE_31), .ZN(n36) );
  INV_X1 U36 ( .A(INSTR_EXE[19]), .ZN(n27) );
  INV_X1 U37 ( .A(INSTR_EXE[16]), .ZN(n26) );
  INV_X1 U38 ( .A(INSTR_EXE[20]), .ZN(n25) );
  INV_X1 U39 ( .A(INSTR_EXE[18]), .ZN(n28) );
  INV_X1 U40 ( .A(INSTR_EXE_31), .ZN(n31) );
  INV_X1 U41 ( .A(INSTR_EXE_30), .ZN(n30) );
  AOI221_X1 U42 ( .B1(INSTR_EXE_30), .B2(n31), .C1(n30), .C2(INSTR_EXE_31), 
        .A(n29), .ZN(n32) );
  NAND3_X1 U43 ( .A1(INSTR_EXE_27), .A2(INSTR_EXE_28), .A3(n32), .ZN(n37) );
  INV_X1 U44 ( .A(n36), .ZN(n38) );
  NAND4_X1 U45 ( .A1(INSTR_EXE_4), .A2(INSTR_EXE_2), .A3(INSTR_EXE_1), .A4(
        INSTR_EXE_3), .ZN(n33) );
  AOI221_X1 U46 ( .B1(n38), .B2(n37), .C1(n36), .C2(n35), .A(INSTR_EXE_26), 
        .ZN(N683) );
  INV_X1 U47 ( .A(\HDU_OUTS[PC_EN] ), .ZN(n39) );
endmodule


module FU ( INSTR_ID, INSTR_EXE, INSTR_MEM, INSTR_WB, .FU_OUTS({
        \FU_OUTS[MUX_RF_OUT1_SEL][2] , \FU_OUTS[MUX_RF_OUT1_SEL][1] , 
        \FU_OUTS[MUX_RF_OUT1_SEL][0] , \FU_OUTS[MUX_RF_OUT2_SEL][2] , 
        \FU_OUTS[MUX_RF_OUT2_SEL][1] , \FU_OUTS[MUX_RF_OUT2_SEL][0] , 
        \FU_OUTS[MUX_DRAM_IN_SEL] }) );
  input [31:0] INSTR_ID;
  input [31:0] INSTR_EXE;
  input [31:0] INSTR_MEM;
  input [31:0] INSTR_WB;
  output \FU_OUTS[MUX_RF_OUT1_SEL][2] , \FU_OUTS[MUX_RF_OUT1_SEL][1] ,
         \FU_OUTS[MUX_RF_OUT1_SEL][0] , \FU_OUTS[MUX_RF_OUT2_SEL][2] ,
         \FU_OUTS[MUX_RF_OUT2_SEL][1] , \FU_OUTS[MUX_RF_OUT2_SEL][0] ,
         \FU_OUTS[MUX_DRAM_IN_SEL] ;
  wire   INSTR_EXE_31, INSTR_EXE_30, INSTR_EXE_29, INSTR_EXE_28, INSTR_EXE_27,
         INSTR_EXE_26, INSTR_MEM_31, INSTR_MEM_30, INSTR_MEM_29, INSTR_MEM_28,
         INSTR_MEM_27, INSTR_MEM_26, INSTR_WB_31, INSTR_WB_30, INSTR_WB_29,
         INSTR_WB_28, INSTR_WB_27, INSTR_WB_26, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159;
  assign INSTR_EXE_31 = INSTR_EXE[31];
  assign INSTR_EXE_30 = INSTR_EXE[30];
  assign INSTR_EXE_29 = INSTR_EXE[29];
  assign INSTR_EXE_28 = INSTR_EXE[28];
  assign INSTR_EXE_27 = INSTR_EXE[27];
  assign INSTR_EXE_26 = INSTR_EXE[26];
  assign INSTR_MEM_31 = INSTR_MEM[31];
  assign INSTR_MEM_30 = INSTR_MEM[30];
  assign INSTR_MEM_29 = INSTR_MEM[29];
  assign INSTR_MEM_28 = INSTR_MEM[28];
  assign INSTR_MEM_27 = INSTR_MEM[27];
  assign INSTR_MEM_26 = INSTR_MEM[26];
  assign INSTR_WB_31 = INSTR_WB[31];
  assign INSTR_WB_30 = INSTR_WB[30];
  assign INSTR_WB_29 = INSTR_WB[29];
  assign INSTR_WB_28 = INSTR_WB[28];
  assign INSTR_WB_27 = INSTR_WB[27];
  assign INSTR_WB_26 = INSTR_WB[26];

  AOI21_X1 U3 ( .B1(n156), .B2(n158), .A(n132), .ZN(
        \FU_OUTS[MUX_RF_OUT2_SEL][1] ) );
  INV_X1 U4 ( .A(n57), .ZN(\FU_OUTS[MUX_RF_OUT1_SEL][1] ) );
  NOR3_X1 U5 ( .A1(n17), .A2(n16), .A3(n15), .ZN(\FU_OUTS[MUX_DRAM_IN_SEL] )
         );
  OAI21_X1 U6 ( .B1(n82), .B2(n81), .A(n80), .ZN(\FU_OUTS[MUX_RF_OUT1_SEL][2] ) );
  AND2_X1 U7 ( .A1(n51), .A2(n1), .ZN(n82) );
  AND3_X1 U8 ( .A1(n22), .A2(n23), .A3(n2), .ZN(n51) );
  INV_X1 U9 ( .A(n9), .ZN(n8) );
  NOR2_X1 U10 ( .A1(n84), .A2(n75), .ZN(n79) );
  INV_X1 U11 ( .A(INSTR_EXE_28), .ZN(n35) );
  INV_X1 U12 ( .A(INSTR_MEM_29), .ZN(n125) );
  NOR4_X2 U13 ( .A1(INSTR_WB_30), .A2(INSTR_WB_29), .A3(INSTR_WB_27), .A4(n58), 
        .ZN(n68) );
  OAI221_X1 U14 ( .B1(n79), .B2(n74), .C1(n79), .C2(n48), .A(n76), .ZN(
        \FU_OUTS[MUX_RF_OUT1_SEL][0] ) );
  INV_X1 U15 ( .A(n43), .ZN(n42) );
  NOR4_X2 U16 ( .A1(INSTR_EXE_26), .A2(INSTR_EXE_27), .A3(INSTR_EXE_30), .A4(
        n30), .ZN(n43) );
  INV_X1 U17 ( .A(n33), .ZN(n30) );
  NOR2_X1 U18 ( .A1(INSTR_EXE_29), .A2(INSTR_EXE_31), .ZN(n33) );
  OR2_X1 U19 ( .A1(INSTR_WB_26), .A2(INSTR_WB_31), .ZN(n58) );
  AOI22_X1 U20 ( .A1(n9), .A2(INSTR_MEM[12]), .B1(INSTR_MEM[17]), .B2(n8), 
        .ZN(n94) );
  AOI22_X1 U21 ( .A1(n9), .A2(INSTR_MEM[14]), .B1(INSTR_MEM[19]), .B2(n8), 
        .ZN(n91) );
  AOI22_X1 U22 ( .A1(n9), .A2(INSTR_MEM[13]), .B1(INSTR_MEM[18]), .B2(n8), 
        .ZN(n97) );
  AOI22_X1 U23 ( .A1(n9), .A2(INSTR_MEM[15]), .B1(INSTR_MEM[20]), .B2(n8), 
        .ZN(n96) );
  NOR2_X2 U24 ( .A1(INSTR_MEM_26), .A2(n54), .ZN(n9) );
  NAND3_X1 U25 ( .A1(n107), .A2(n10), .A3(n52), .ZN(n54) );
  OAI21_X1 U26 ( .B1(INSTR_MEM_28), .B2(n125), .A(n25), .ZN(n52) );
  AOI21_X1 U27 ( .B1(INSTR_MEM_31), .B2(INSTR_MEM_30), .A(n104), .ZN(n25) );
  INV_X1 U28 ( .A(INSTR_MEM_27), .ZN(n104) );
  OR3_X1 U29 ( .A1(n75), .A2(n19), .A3(n87), .ZN(n74) );
  INV_X1 U30 ( .A(INSTR_MEM_30), .ZN(n10) );
  NOR2_X1 U31 ( .A1(INSTR_MEM_31), .A2(INSTR_MEM_29), .ZN(n107) );
  OR4_X1 U32 ( .A1(INSTR_ID[21]), .A2(INSTR_ID[22]), .A3(INSTR_ID[25]), .A4(
        INSTR_ID[23]), .ZN(n24) );
  NOR3_X1 U33 ( .A1(n55), .A2(n56), .A3(n123), .ZN(n1) );
  INV_X1 U34 ( .A(n54), .ZN(n5) );
  NOR2_X1 U35 ( .A1(n53), .A2(n52), .ZN(n4) );
  XNOR2_X1 U36 ( .A(n93), .B(n3), .ZN(n2) );
  INV_X1 U37 ( .A(INSTR_ID[21]), .ZN(n3) );
  MUX2_X1 U38 ( .A(n4), .B(n5), .S(INSTR_MEM_28), .Z(n55) );
  AOI22_X1 U39 ( .A1(INSTR_EXE[18]), .A2(n97), .B1(INSTR_EXE[19]), .B2(n91), 
        .ZN(n6) );
  OAI221_X1 U40 ( .B1(INSTR_EXE[18]), .B2(n97), .C1(INSTR_EXE[19]), .C2(n91), 
        .A(n6), .ZN(n17) );
  AOI22_X1 U41 ( .A1(n9), .A2(INSTR_MEM[11]), .B1(INSTR_MEM[16]), .B2(n8), 
        .ZN(n93) );
  AOI22_X1 U42 ( .A1(INSTR_EXE[20]), .A2(n96), .B1(INSTR_EXE[16]), .B2(n93), 
        .ZN(n7) );
  OAI221_X1 U43 ( .B1(INSTR_EXE[20]), .B2(n96), .C1(INSTR_EXE[16]), .C2(n93), 
        .A(n7), .ZN(n16) );
  INV_X1 U44 ( .A(INSTR_MEM_28), .ZN(n122) );
  AOI21_X1 U45 ( .B1(n122), .B2(INSTR_MEM_26), .A(n104), .ZN(n87) );
  NAND2_X1 U46 ( .A1(n10), .A2(INSTR_MEM_31), .ZN(n49) );
  INV_X1 U47 ( .A(n49), .ZN(n53) );
  NAND2_X1 U48 ( .A1(n53), .A2(n125), .ZN(n86) );
  NAND2_X1 U49 ( .A1(INSTR_MEM_27), .A2(INSTR_MEM_28), .ZN(n11) );
  NOR3_X1 U50 ( .A1(INSTR_MEM_31), .A2(INSTR_MEM_30), .A3(n125), .ZN(n85) );
  NAND2_X1 U51 ( .A1(INSTR_MEM_26), .A2(n85), .ZN(n27) );
  OAI22_X1 U52 ( .A1(n87), .A2(n86), .B1(n11), .B2(n27), .ZN(n14) );
  INV_X1 U53 ( .A(n91), .ZN(n89) );
  NOR4_X1 U54 ( .A1(INSTR_EXE[16]), .A2(INSTR_EXE[20]), .A3(INSTR_EXE[18]), 
        .A4(n89), .ZN(n12) );
  OAI21_X1 U55 ( .B1(INSTR_EXE[17]), .B2(n12), .A(n94), .ZN(n13) );
  OAI211_X1 U56 ( .C1(INSTR_EXE[17]), .C2(n94), .A(n14), .B(n13), .ZN(n15) );
  NAND4_X1 U57 ( .A1(INSTR_EXE_27), .A2(n33), .A3(INSTR_EXE_26), .A4(n35), 
        .ZN(n84) );
  AND2_X1 U58 ( .A1(INSTR_ID[25]), .A2(INSTR_ID[23]), .ZN(n18) );
  NAND4_X1 U59 ( .A1(INSTR_ID[24]), .A2(INSTR_ID[21]), .A3(INSTR_ID[22]), .A4(
        n18), .ZN(n75) );
  NOR4_X1 U60 ( .A1(INSTR_MEM_31), .A2(INSTR_MEM_28), .A3(INSTR_MEM_29), .A4(
        n104), .ZN(n126) );
  INV_X1 U61 ( .A(n126), .ZN(n19) );
  OAI22_X1 U62 ( .A1(INSTR_ID[24]), .A2(n91), .B1(INSTR_ID[22]), .B2(n94), 
        .ZN(n20) );
  AOI221_X1 U63 ( .B1(INSTR_ID[24]), .B2(n91), .C1(n94), .C2(INSTR_ID[22]), 
        .A(n20), .ZN(n23) );
  OAI22_X1 U64 ( .A1(INSTR_ID[25]), .A2(n96), .B1(INSTR_ID[23]), .B2(n97), 
        .ZN(n21) );
  AOI221_X1 U65 ( .B1(INSTR_ID[25]), .B2(n96), .C1(n97), .C2(INSTR_ID[23]), 
        .A(n21), .ZN(n22) );
  NOR2_X1 U66 ( .A1(n24), .A2(INSTR_ID[24]), .ZN(n56) );
  INV_X1 U67 ( .A(n56), .ZN(n63) );
  INV_X1 U68 ( .A(INSTR_MEM_26), .ZN(n103) );
  OAI21_X1 U69 ( .B1(n103), .B2(INSTR_MEM_28), .A(n25), .ZN(n26) );
  INV_X1 U70 ( .A(n26), .ZN(n28) );
  OAI22_X1 U71 ( .A1(n28), .A2(n86), .B1(n52), .B2(n27), .ZN(n29) );
  NAND3_X1 U72 ( .A1(n51), .A2(n63), .A3(n29), .ZN(n48) );
  AOI22_X1 U73 ( .A1(n43), .A2(INSTR_EXE[12]), .B1(INSTR_EXE[17]), .B2(n42), 
        .ZN(n110) );
  AOI22_X1 U74 ( .A1(n43), .A2(INSTR_EXE[15]), .B1(INSTR_EXE[20]), .B2(n42), 
        .ZN(n114) );
  OAI22_X1 U75 ( .A1(n110), .A2(INSTR_ID[22]), .B1(n114), .B2(INSTR_ID[25]), 
        .ZN(n31) );
  AOI221_X1 U76 ( .B1(n110), .B2(INSTR_ID[22]), .C1(INSTR_ID[25]), .C2(n114), 
        .A(n31), .ZN(n47) );
  AOI22_X1 U77 ( .A1(n43), .A2(INSTR_EXE[13]), .B1(INSTR_EXE[18]), .B2(n42), 
        .ZN(n109) );
  INV_X1 U78 ( .A(INSTR_EXE_30), .ZN(n32) );
  NAND4_X1 U79 ( .A1(INSTR_EXE_31), .A2(INSTR_EXE_29), .A3(n32), .A4(n35), 
        .ZN(n37) );
  NOR2_X1 U80 ( .A1(INSTR_EXE_27), .A2(n37), .ZN(n40) );
  INV_X1 U81 ( .A(INSTR_EXE_26), .ZN(n38) );
  NOR2_X1 U82 ( .A1(INSTR_EXE_27), .A2(INSTR_EXE_30), .ZN(n34) );
  OAI221_X1 U83 ( .B1(INSTR_EXE_28), .B2(INSTR_EXE_27), .C1(n35), .C2(n34), 
        .A(n33), .ZN(n36) );
  OAI21_X1 U84 ( .B1(n38), .B2(n37), .A(n36), .ZN(n39) );
  NOR2_X1 U85 ( .A1(n40), .A2(n39), .ZN(n121) );
  OAI211_X1 U86 ( .C1(n109), .C2(INSTR_ID[23]), .A(n121), .B(n63), .ZN(n41) );
  AOI21_X1 U87 ( .B1(n109), .B2(INSTR_ID[23]), .A(n41), .ZN(n46) );
  AOI22_X1 U88 ( .A1(n43), .A2(INSTR_EXE[14]), .B1(INSTR_EXE[19]), .B2(n42), 
        .ZN(n117) );
  AOI22_X1 U89 ( .A1(n43), .A2(INSTR_EXE[11]), .B1(INSTR_EXE[16]), .B2(n42), 
        .ZN(n116) );
  OAI22_X1 U90 ( .A1(n117), .A2(INSTR_ID[24]), .B1(n116), .B2(INSTR_ID[21]), 
        .ZN(n44) );
  AOI221_X1 U91 ( .B1(n117), .B2(INSTR_ID[24]), .C1(INSTR_ID[21]), .C2(n116), 
        .A(n44), .ZN(n45) );
  NAND3_X1 U92 ( .A1(n47), .A2(n46), .A3(n45), .ZN(n76) );
  NAND2_X1 U93 ( .A1(INSTR_MEM_29), .A2(n122), .ZN(n50) );
  AOI211_X1 U94 ( .C1(INSTR_MEM_27), .C2(n103), .A(n50), .B(n49), .ZN(n123) );
  OAI21_X1 U95 ( .B1(n79), .B2(n82), .A(n76), .ZN(n57) );
  INV_X1 U96 ( .A(n68), .ZN(n67) );
  AOI22_X1 U97 ( .A1(n68), .A2(INSTR_WB[15]), .B1(INSTR_WB[20]), .B2(n67), 
        .ZN(n146) );
  AOI22_X1 U98 ( .A1(n68), .A2(INSTR_WB[11]), .B1(INSTR_WB[16]), .B2(n67), 
        .ZN(n143) );
  AOI22_X1 U99 ( .A1(INSTR_ID[25]), .A2(n146), .B1(INSTR_ID[21]), .B2(n143), 
        .ZN(n59) );
  OAI221_X1 U100 ( .B1(INSTR_ID[25]), .B2(n146), .C1(INSTR_ID[21]), .C2(n143), 
        .A(n59), .ZN(n72) );
  AOI22_X1 U101 ( .A1(n68), .A2(INSTR_WB[12]), .B1(INSTR_WB[17]), .B2(n67), 
        .ZN(n145) );
  INV_X1 U102 ( .A(INSTR_WB_27), .ZN(n138) );
  NOR4_X1 U103 ( .A1(INSTR_WB_29), .A2(INSTR_WB_28), .A3(INSTR_WB_31), .A4(
        n138), .ZN(n73) );
  INV_X1 U104 ( .A(INSTR_WB_28), .ZN(n60) );
  NOR3_X1 U105 ( .A1(INSTR_WB_30), .A2(INSTR_WB_29), .A3(n60), .ZN(n139) );
  NAND2_X1 U106 ( .A1(n139), .A2(n138), .ZN(n64) );
  INV_X1 U107 ( .A(INSTR_WB_29), .ZN(n61) );
  NOR3_X1 U108 ( .A1(INSTR_WB_30), .A2(INSTR_WB_28), .A3(n61), .ZN(n62) );
  OAI211_X1 U109 ( .C1(INSTR_WB_26), .C2(n138), .A(INSTR_WB_31), .B(n62), .ZN(
        n147) );
  OAI211_X1 U110 ( .C1(INSTR_WB_31), .C2(n64), .A(n63), .B(n147), .ZN(n65) );
  AOI211_X1 U111 ( .C1(n145), .C2(INSTR_ID[22]), .A(n73), .B(n65), .ZN(n66) );
  OAI21_X1 U112 ( .B1(n145), .B2(INSTR_ID[22]), .A(n66), .ZN(n71) );
  AOI22_X1 U113 ( .A1(n68), .A2(INSTR_WB[13]), .B1(INSTR_WB[18]), .B2(n67), 
        .ZN(n135) );
  AOI22_X1 U114 ( .A1(n68), .A2(INSTR_WB[14]), .B1(INSTR_WB[19]), .B2(n67), 
        .ZN(n134) );
  AOI22_X1 U115 ( .A1(INSTR_ID[23]), .A2(n135), .B1(INSTR_ID[24]), .B2(n134), 
        .ZN(n69) );
  OAI221_X1 U116 ( .B1(INSTR_ID[23]), .B2(n135), .C1(INSTR_ID[24]), .C2(n134), 
        .A(n69), .ZN(n70) );
  NOR3_X1 U117 ( .A1(n72), .A2(n71), .A3(n70), .ZN(n78) );
  NAND2_X1 U118 ( .A1(INSTR_WB_26), .A2(n73), .ZN(n153) );
  OAI21_X1 U119 ( .B1(n75), .B2(n153), .A(n74), .ZN(n77) );
  OAI21_X1 U120 ( .B1(n78), .B2(n77), .A(n76), .ZN(n81) );
  INV_X1 U121 ( .A(n79), .ZN(n80) );
  AND2_X1 U122 ( .A1(INSTR_ID[17]), .A2(INSTR_ID[20]), .ZN(n83) );
  NAND4_X1 U123 ( .A1(INSTR_ID[19]), .A2(INSTR_ID[16]), .A3(INSTR_ID[18]), 
        .A4(n83), .ZN(n154) );
  NOR2_X1 U124 ( .A1(n84), .A2(n154), .ZN(n131) );
  AND4_X1 U125 ( .A1(INSTR_MEM_27), .A2(INSTR_MEM_26), .A3(INSTR_MEM_28), .A4(
        n85), .ZN(n102) );
  NOR3_X1 U126 ( .A1(n87), .A2(n126), .A3(n86), .ZN(n101) );
  INV_X1 U127 ( .A(INSTR_ID[19]), .ZN(n90) );
  OR4_X1 U128 ( .A1(INSTR_ID[19]), .A2(INSTR_ID[18]), .A3(INSTR_ID[17]), .A4(
        INSTR_ID[20]), .ZN(n88) );
  NOR2_X1 U129 ( .A1(n88), .A2(INSTR_ID[16]), .ZN(n111) );
  INV_X1 U130 ( .A(n111), .ZN(n140) );
  OAI221_X1 U131 ( .B1(INSTR_ID[19]), .B2(n91), .C1(n90), .C2(n89), .A(n140), 
        .ZN(n100) );
  AOI22_X1 U132 ( .A1(n94), .A2(INSTR_ID[17]), .B1(n93), .B2(INSTR_ID[16]), 
        .ZN(n92) );
  OAI221_X1 U133 ( .B1(n94), .B2(INSTR_ID[17]), .C1(n93), .C2(INSTR_ID[16]), 
        .A(n92), .ZN(n99) );
  AOI22_X1 U134 ( .A1(n97), .A2(INSTR_ID[18]), .B1(n96), .B2(INSTR_ID[20]), 
        .ZN(n95) );
  OAI221_X1 U135 ( .B1(n97), .B2(INSTR_ID[18]), .C1(n96), .C2(INSTR_ID[20]), 
        .A(n95), .ZN(n98) );
  NOR3_X1 U136 ( .A1(n100), .A2(n99), .A3(n98), .ZN(n130) );
  OAI21_X1 U137 ( .B1(n102), .B2(n101), .A(n130), .ZN(n127) );
  INV_X1 U138 ( .A(n154), .ZN(n106) );
  NOR2_X1 U139 ( .A1(n104), .A2(n103), .ZN(n105) );
  NAND4_X1 U140 ( .A1(n107), .A2(n106), .A3(n105), .A4(n122), .ZN(n152) );
  OAI22_X1 U141 ( .A1(n110), .A2(INSTR_ID[17]), .B1(INSTR_ID[18]), .B2(n109), 
        .ZN(n108) );
  AOI221_X1 U142 ( .B1(n110), .B2(INSTR_ID[17]), .C1(n109), .C2(INSTR_ID[18]), 
        .A(n108), .ZN(n120) );
  INV_X1 U143 ( .A(INSTR_ID[20]), .ZN(n113) );
  INV_X1 U144 ( .A(n114), .ZN(n112) );
  AOI221_X1 U145 ( .B1(INSTR_ID[20]), .B2(n114), .C1(n113), .C2(n112), .A(n111), .ZN(n119) );
  OAI22_X1 U146 ( .A1(n117), .A2(INSTR_ID[19]), .B1(n116), .B2(INSTR_ID[16]), 
        .ZN(n115) );
  AOI221_X1 U147 ( .B1(n117), .B2(INSTR_ID[19]), .C1(INSTR_ID[16]), .C2(n116), 
        .A(n115), .ZN(n118) );
  NAND4_X1 U148 ( .A1(n121), .A2(n120), .A3(n119), .A4(n118), .ZN(n157) );
  OAI221_X1 U149 ( .B1(n131), .B2(n127), .C1(n131), .C2(n152), .A(n157), .ZN(
        \FU_OUTS[MUX_RF_OUT2_SEL][0] ) );
  NOR3_X1 U150 ( .A1(INSTR_MEM_27), .A2(INSTR_MEM_30), .A3(n122), .ZN(n124) );
  AOI221_X1 U151 ( .B1(n126), .B2(n125), .C1(n124), .C2(n125), .A(n123), .ZN(
        n129) );
  INV_X1 U152 ( .A(n127), .ZN(n128) );
  AOI21_X1 U153 ( .B1(n130), .B2(n129), .A(n128), .ZN(n156) );
  INV_X1 U154 ( .A(n131), .ZN(n158) );
  INV_X1 U155 ( .A(n157), .ZN(n132) );
  OAI22_X1 U156 ( .A1(n135), .A2(INSTR_ID[18]), .B1(INSTR_ID[19]), .B2(n134), 
        .ZN(n133) );
  AOI221_X1 U157 ( .B1(n135), .B2(INSTR_ID[18]), .C1(n134), .C2(INSTR_ID[19]), 
        .A(n133), .ZN(n150) );
  NOR2_X1 U158 ( .A1(INSTR_WB_29), .A2(INSTR_WB_28), .ZN(n137) );
  INV_X1 U159 ( .A(INSTR_WB_31), .ZN(n136) );
  OAI221_X1 U160 ( .B1(INSTR_WB_27), .B2(n139), .C1(n138), .C2(n137), .A(n136), 
        .ZN(n141) );
  OAI211_X1 U161 ( .C1(n143), .C2(INSTR_ID[16]), .A(n141), .B(n140), .ZN(n142)
         );
  AOI21_X1 U162 ( .B1(n143), .B2(INSTR_ID[16]), .A(n142), .ZN(n149) );
  OAI22_X1 U163 ( .A1(n146), .A2(INSTR_ID[20]), .B1(INSTR_ID[17]), .B2(n145), 
        .ZN(n144) );
  AOI221_X1 U164 ( .B1(n146), .B2(INSTR_ID[20]), .C1(n145), .C2(INSTR_ID[17]), 
        .A(n144), .ZN(n148) );
  NAND4_X1 U165 ( .A1(n150), .A2(n149), .A3(n148), .A4(n147), .ZN(n151) );
  OAI211_X1 U166 ( .C1(n154), .C2(n153), .A(n152), .B(n151), .ZN(n155) );
  NAND3_X1 U167 ( .A1(n157), .A2(n156), .A3(n155), .ZN(n159) );
  NAND2_X1 U168 ( .A1(n159), .A2(n158), .ZN(\FU_OUTS[MUX_RF_OUT2_SEL][2] ) );
endmodule


module CU ( INSTR_ID, .CU_OUTS({\CU_OUTS[ID][MUX_BRANCH_SEL] , 
        \CU_OUTS[ID][MUX_IMM_EXT_SEL] , \CU_OUTS[ID][MUX_RF_WR_ADDR_SEL][1] , 
        \CU_OUTS[ID][MUX_RF_WR_ADDR_SEL][0] , \CU_OUTS[ID][BRANCH_COND][1] , 
        \CU_OUTS[ID][BRANCH_COND][0] , \CU_OUTS[EXE][MULT_EN] , 
        \CU_OUTS[EXE][MUX_MULT_SEL] , \CU_OUTS[EXE][MUX_ALU_IN2_SEL] , 
        \CU_OUTS[EXE][ALU_OP][4] , \CU_OUTS[EXE][ALU_OP][3] , 
        \CU_OUTS[EXE][ALU_OP][2] , \CU_OUTS[EXE][ALU_OP][1] , 
        \CU_OUTS[EXE][ALU_OP][0] , \CU_OUTS[MEM][DRAM_WR_EN][1] , 
        \CU_OUTS[MEM][DRAM_WR_EN][0] , \CU_OUTS[MEM][MUX_DRAM_OUT_EXT_SEL][2] , 
        \CU_OUTS[MEM][MUX_DRAM_OUT_EXT_SEL][1] , 
        \CU_OUTS[MEM][MUX_DRAM_OUT_EXT_SEL][0] , \CU_OUTS[WB][MUX_WB_SEL][1] , 
        \CU_OUTS[WB][MUX_WB_SEL][0] , \CU_OUTS[WB][RF_WR_EN] }) );
  input [31:0] INSTR_ID;
  output \CU_OUTS[ID][MUX_BRANCH_SEL] , \CU_OUTS[ID][MUX_IMM_EXT_SEL] ,
         \CU_OUTS[ID][MUX_RF_WR_ADDR_SEL][1] ,
         \CU_OUTS[ID][MUX_RF_WR_ADDR_SEL][0] , \CU_OUTS[ID][BRANCH_COND][1] ,
         \CU_OUTS[ID][BRANCH_COND][0] , \CU_OUTS[EXE][MULT_EN] ,
         \CU_OUTS[EXE][MUX_MULT_SEL] , \CU_OUTS[EXE][MUX_ALU_IN2_SEL] ,
         \CU_OUTS[EXE][ALU_OP][4] , \CU_OUTS[EXE][ALU_OP][3] ,
         \CU_OUTS[EXE][ALU_OP][2] , \CU_OUTS[EXE][ALU_OP][1] ,
         \CU_OUTS[EXE][ALU_OP][0] , \CU_OUTS[MEM][DRAM_WR_EN][1] ,
         \CU_OUTS[MEM][DRAM_WR_EN][0] ,
         \CU_OUTS[MEM][MUX_DRAM_OUT_EXT_SEL][2] ,
         \CU_OUTS[MEM][MUX_DRAM_OUT_EXT_SEL][1] ,
         \CU_OUTS[MEM][MUX_DRAM_OUT_EXT_SEL][0] , \CU_OUTS[WB][MUX_WB_SEL][1] ,
         \CU_OUTS[WB][MUX_WB_SEL][0] , \CU_OUTS[WB][RF_WR_EN] ;
  wire   INSTR_ID_5, INSTR_ID_4, INSTR_ID_3, INSTR_ID_2, INSTR_ID_1,
         INSTR_ID_0, \CU_OUTS[ID][MUX_IMM_EXT_SEL] , \INSTR_ID[27] ,
         \INSTR_ID[28] , n96, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95;
  assign INSTR_ID_5 = INSTR_ID[5];
  assign INSTR_ID_4 = INSTR_ID[4];
  assign INSTR_ID_3 = INSTR_ID[3];
  assign INSTR_ID_2 = INSTR_ID[2];
  assign INSTR_ID_1 = INSTR_ID[1];
  assign INSTR_ID_0 = INSTR_ID[0];
  assign \CU_OUTS[ID][MUX_RF_WR_ADDR_SEL][1]  = \CU_OUTS[ID][MUX_IMM_EXT_SEL] ;
  assign \CU_OUTS[MEM][MUX_DRAM_OUT_EXT_SEL][2]  = \INSTR_ID[27] ;
  assign \INSTR_ID[27]  = INSTR_ID[27];
  assign \CU_OUTS[MEM][MUX_DRAM_OUT_EXT_SEL][0]  = \INSTR_ID[28] ;
  assign \INSTR_ID[28]  = INSTR_ID[28];

  XOR2_X1 U3 ( .A(\INSTR_ID[28] ), .B(\INSTR_ID[27] ), .Z(n18) );
  INV_X1 U4 ( .A(INSTR_ID_1), .ZN(n1) );
  NAND4_X1 U5 ( .A1(INSTR_ID_5), .A2(INSTR_ID_3), .A3(n14), .A4(INSTR_ID_2), 
        .ZN(n2) );
  OAI21_X1 U6 ( .B1(n1), .B2(n2), .A(n12), .ZN(n35) );
  OR2_X1 U7 ( .A1(n52), .A2(INSTR_ID[30]), .ZN(n54) );
  INV_X1 U8 ( .A(INSTR_ID[29]), .ZN(n65) );
  INV_X1 U9 ( .A(INSTR_ID[31]), .ZN(n50) );
  INV_X1 U10 ( .A(INSTR_ID[26]), .ZN(n73) );
  NOR3_X4 U11 ( .A1(\INSTR_ID[28] ), .A2(\CU_OUTS[ID][MUX_RF_WR_ADDR_SEL][0] ), 
        .A3(n52), .ZN(\CU_OUTS[ID][MUX_IMM_EXT_SEL] ) );
  NAND2_X1 U12 ( .A1(n50), .A2(n65), .ZN(n52) );
  INV_X1 U13 ( .A(\INSTR_ID[28] ), .ZN(n63) );
  NOR4_X2 U14 ( .A1(\INSTR_ID[27] ), .A2(INSTR_ID[26]), .A3(\INSTR_ID[28] ), 
        .A4(n54), .ZN(\CU_OUTS[ID][MUX_RF_WR_ADDR_SEL][0] ) );
  NOR2_X1 U15 ( .A1(\INSTR_ID[27] ), .A2(n73), .ZN(
        \CU_OUTS[MEM][MUX_DRAM_OUT_EXT_SEL][1] ) );
  NOR2_X1 U16 ( .A1(INSTR_ID[30]), .A2(n50), .ZN(\CU_OUTS[WB][MUX_WB_SEL][0] )
         );
  INV_X1 U17 ( .A(\CU_OUTS[ID][MUX_RF_WR_ADDR_SEL][0] ), .ZN(n96) );
  INV_X1 U18 ( .A(INSTR_ID_5), .ZN(n3) );
  INV_X1 U19 ( .A(INSTR_ID_3), .ZN(n4) );
  AOI21_X1 U20 ( .B1(INSTR_ID_2), .B2(n3), .A(n4), .ZN(n16) );
  INV_X1 U21 ( .A(INSTR_ID_4), .ZN(n14) );
  AOI21_X1 U22 ( .B1(INSTR_ID_5), .B2(n4), .A(n14), .ZN(n9) );
  AOI211_X1 U23 ( .C1(INSTR_ID_0), .C2(n16), .A(INSTR_ID_1), .B(n9), .ZN(n11)
         );
  NOR2_X1 U24 ( .A1(INSTR_ID_4), .A2(INSTR_ID_3), .ZN(n7) );
  AOI21_X1 U25 ( .B1(INSTR_ID_4), .B2(n4), .A(n3), .ZN(n12) );
  OAI221_X1 U26 ( .B1(INSTR_ID_4), .B2(INSTR_ID_5), .C1(n14), .C2(INSTR_ID_3), 
        .A(INSTR_ID_2), .ZN(n5) );
  AOI21_X1 U27 ( .B1(INSTR_ID_1), .B2(n12), .A(n5), .ZN(n6) );
  AOI21_X1 U28 ( .B1(n7), .B2(INSTR_ID_2), .A(n6), .ZN(n85) );
  INV_X1 U29 ( .A(n9), .ZN(n82) );
  NAND4_X1 U30 ( .A1(INSTR_ID_5), .A2(INSTR_ID_4), .A3(INSTR_ID_3), .A4(
        INSTR_ID_2), .ZN(n8) );
  NAND2_X1 U31 ( .A1(INSTR_ID_1), .A2(n8), .ZN(n84) );
  NAND2_X1 U32 ( .A1(n85), .A2(n84), .ZN(n13) );
  NAND2_X1 U33 ( .A1(n16), .A2(n13), .ZN(n59) );
  NOR3_X1 U34 ( .A1(n9), .A2(n85), .A3(n16), .ZN(n38) );
  INV_X1 U35 ( .A(INSTR_ID_0), .ZN(n91) );
  NAND2_X1 U36 ( .A1(n38), .A2(n91), .ZN(n62) );
  OAI22_X1 U37 ( .A1(n82), .A2(n59), .B1(n84), .B2(n62), .ZN(n10) );
  AOI221_X1 U38 ( .B1(INSTR_ID_0), .B2(n11), .C1(n85), .C2(n11), .A(n10), .ZN(
        n25) );
  NOR2_X1 U39 ( .A1(n96), .A2(n35), .ZN(n83) );
  INV_X1 U40 ( .A(n83), .ZN(n60) );
  INV_X1 U41 ( .A(n13), .ZN(n15) );
  NAND3_X1 U42 ( .A1(n16), .A2(n15), .A3(n14), .ZN(n61) );
  INV_X1 U43 ( .A(n84), .ZN(n34) );
  NAND2_X1 U44 ( .A1(n34), .A2(n38), .ZN(n89) );
  NAND2_X1 U45 ( .A1(\CU_OUTS[ID][MUX_RF_WR_ADDR_SEL][0] ), .A2(n35), .ZN(n88)
         );
  AOI21_X1 U46 ( .B1(n61), .B2(n89), .A(n88), .ZN(n42) );
  INV_X1 U47 ( .A(\INSTR_ID[27] ), .ZN(n70) );
  INV_X1 U48 ( .A(INSTR_ID[30]), .ZN(n64) );
  NOR3_X1 U49 ( .A1(INSTR_ID[31]), .A2(n64), .A3(n63), .ZN(n75) );
  OAI211_X1 U50 ( .C1(INSTR_ID[26]), .C2(n70), .A(n75), .B(n65), .ZN(n17) );
  NAND3_X1 U51 ( .A1(INSTR_ID[29]), .A2(INSTR_ID[30]), .A3(n18), .ZN(n94) );
  OAI22_X1 U52 ( .A1(\CU_OUTS[MEM][MUX_DRAM_OUT_EXT_SEL][1] ), .A2(n17), .B1(
        n50), .B2(n94), .ZN(n23) );
  NOR3_X1 U53 ( .A1(\INSTR_ID[27] ), .A2(\INSTR_ID[28] ), .A3(n65), .ZN(n56)
         );
  NOR2_X1 U54 ( .A1(INSTR_ID[31]), .A2(n65), .ZN(n71) );
  OAI221_X1 U55 ( .B1(n56), .B2(n71), .C1(n56), .C2(
        \CU_OUTS[MEM][MUX_DRAM_OUT_EXT_SEL][1] ), .A(n64), .ZN(n21) );
  NAND3_X1 U56 ( .A1(INSTR_ID[26]), .A2(\CU_OUTS[WB][MUX_WB_SEL][0] ), .A3(n63), .ZN(n55) );
  NAND3_X1 U57 ( .A1(\CU_OUTS[WB][MUX_WB_SEL][0] ), .A2(n65), .A3(n70), .ZN(
        n68) );
  INV_X1 U58 ( .A(n18), .ZN(n19) );
  NAND3_X1 U59 ( .A1(n71), .A2(n73), .A3(n19), .ZN(n20) );
  NAND4_X1 U60 ( .A1(n21), .A2(n55), .A3(n68), .A4(n20), .ZN(n22) );
  AOI211_X1 U61 ( .C1(INSTR_ID_0), .C2(n42), .A(n23), .B(n22), .ZN(n24) );
  OR3_X1 U62 ( .A1(n88), .A2(n62), .A3(n34), .ZN(n30) );
  OAI211_X1 U63 ( .C1(n25), .C2(n60), .A(n24), .B(n30), .ZN(
        \CU_OUTS[EXE][ALU_OP][0] ) );
  NOR2_X1 U64 ( .A1(\INSTR_ID[27] ), .A2(n63), .ZN(n32) );
  INV_X1 U65 ( .A(n32), .ZN(n53) );
  NOR4_X1 U66 ( .A1(INSTR_ID[26]), .A2(n64), .A3(n52), .A4(n53), .ZN(n29) );
  NAND3_X1 U67 ( .A1(INSTR_ID[29]), .A2(INSTR_ID[30]), .A3(\INSTR_ID[27] ), 
        .ZN(n47) );
  NOR2_X1 U68 ( .A1(\INSTR_ID[28] ), .A2(n47), .ZN(n44) );
  OAI211_X1 U69 ( .C1(n91), .C2(n85), .A(n34), .B(n83), .ZN(n26) );
  INV_X1 U70 ( .A(n26), .ZN(n28) );
  OAI21_X1 U71 ( .B1(n73), .B2(n63), .A(n71), .ZN(n76) );
  OAI22_X1 U72 ( .A1(INSTR_ID[31]), .A2(n47), .B1(n76), .B2(n70), .ZN(n27) );
  NOR4_X1 U73 ( .A1(n29), .A2(n44), .A3(n28), .A4(n27), .ZN(n31) );
  OAI211_X1 U74 ( .C1(n88), .C2(n61), .A(n31), .B(n30), .ZN(
        \CU_OUTS[EXE][ALU_OP][1] ) );
  NOR2_X1 U75 ( .A1(INSTR_ID[26]), .A2(n52), .ZN(n33) );
  OAI221_X1 U76 ( .B1(INSTR_ID[30]), .B2(n71), .C1(n64), .C2(n33), .A(n32), 
        .ZN(n40) );
  AOI211_X1 U77 ( .C1(INSTR_ID_0), .C2(n35), .A(n34), .B(n96), .ZN(n37) );
  NOR3_X1 U78 ( .A1(n91), .A2(n60), .A3(n59), .ZN(n43) );
  INV_X1 U79 ( .A(n56), .ZN(n36) );
  NAND2_X1 U80 ( .A1(INSTR_ID[30]), .A2(n50), .ZN(n67) );
  OAI22_X1 U81 ( .A1(n60), .A2(n61), .B1(n36), .B2(n67), .ZN(n90) );
  AOI211_X1 U82 ( .C1(n38), .C2(n37), .A(n43), .B(n90), .ZN(n39) );
  OAI211_X1 U83 ( .C1(n73), .C2(n94), .A(n40), .B(n39), .ZN(
        \CU_OUTS[EXE][ALU_OP][2] ) );
  NAND2_X1 U84 ( .A1(INSTR_ID[29]), .A2(INSTR_ID[30]), .ZN(n41) );
  NOR2_X1 U85 ( .A1(n63), .A2(n41), .ZN(n74) );
  AOI22_X1 U86 ( .A1(\INSTR_ID[27] ), .A2(n75), .B1(
        \CU_OUTS[MEM][MUX_DRAM_OUT_EXT_SEL][1] ), .B2(n74), .ZN(n46) );
  AOI211_X1 U87 ( .C1(INSTR_ID[26]), .C2(n44), .A(n43), .B(n42), .ZN(n45) );
  NAND2_X1 U88 ( .A1(n46), .A2(n45), .ZN(\CU_OUTS[EXE][ALU_OP][3] ) );
  OR2_X1 U89 ( .A1(n82), .A2(n88), .ZN(n49) );
  NOR4_X1 U90 ( .A1(n85), .A2(INSTR_ID_0), .A3(n84), .A4(n49), .ZN(n80) );
  NOR4_X1 U91 ( .A1(INSTR_ID[26]), .A2(n50), .A3(n63), .A4(n47), .ZN(n48) );
  OR2_X1 U92 ( .A1(n80), .A2(n48), .ZN(\CU_OUTS[EXE][MULT_EN] ) );
  NAND2_X1 U93 ( .A1(\INSTR_ID[27] ), .A2(\INSTR_ID[28] ), .ZN(n51) );
  OAI21_X1 U94 ( .B1(n51), .B2(n50), .A(n49), .ZN(\CU_OUTS[EXE][MUX_MULT_SEL] ) );
  NOR2_X1 U95 ( .A1(n54), .A2(n53), .ZN(\CU_OUTS[ID][BRANCH_COND][1] ) );
  OAI21_X1 U96 ( .B1(INSTR_ID[30]), .B2(\CU_OUTS[ID][MUX_RF_WR_ADDR_SEL][0] ), 
        .A(n73), .ZN(\CU_OUTS[ID][MUX_BRANCH_SEL] ) );
  NOR2_X1 U97 ( .A1(n65), .A2(n55), .ZN(\CU_OUTS[MEM][DRAM_WR_EN][1] ) );
  INV_X1 U98 ( .A(\CU_OUTS[MEM][DRAM_WR_EN][1] ), .ZN(n58) );
  NAND3_X1 U99 ( .A1(n56), .A2(\CU_OUTS[WB][MUX_WB_SEL][0] ), .A3(n73), .ZN(
        n57) );
  OAI21_X1 U100 ( .B1(n70), .B2(n58), .A(n57), .ZN(
        \CU_OUTS[MEM][DRAM_WR_EN][0] ) );
  OAI211_X1 U101 ( .C1(INSTR_ID[31]), .C2(n63), .A(n96), .B(n65), .ZN(
        \CU_OUTS[WB][MUX_WB_SEL][1] ) );
  NOR2_X1 U102 ( .A1(n60), .A2(n59), .ZN(n92) );
  AOI21_X1 U103 ( .B1(n62), .B2(n61), .A(n96), .ZN(n81) );
  NAND3_X1 U104 ( .A1(n65), .A2(n64), .A3(n63), .ZN(n66) );
  AOI21_X1 U105 ( .B1(n67), .B2(n66), .A(n73), .ZN(n72) );
  INV_X1 U106 ( .A(n68), .ZN(n69) );
  AOI221_X1 U107 ( .B1(n72), .B2(\INSTR_ID[27] ), .C1(n71), .C2(n70), .A(n69), 
        .ZN(n78) );
  OAI21_X1 U108 ( .B1(n75), .B2(n74), .A(n73), .ZN(n77) );
  NAND4_X1 U109 ( .A1(n78), .A2(n94), .A3(n77), .A4(n76), .ZN(n79) );
  NOR4_X1 U110 ( .A1(n92), .A2(n81), .A3(n80), .A4(n79), .ZN(n87) );
  OAI211_X1 U111 ( .C1(n85), .C2(n84), .A(n83), .B(n82), .ZN(n86) );
  OAI211_X1 U112 ( .C1(n89), .C2(n88), .A(n87), .B(n86), .ZN(
        \CU_OUTS[WB][RF_WR_EN] ) );
  AOI21_X1 U113 ( .B1(n92), .B2(n91), .A(n90), .ZN(n93) );
  OAI21_X1 U114 ( .B1(INSTR_ID[26]), .B2(n94), .A(n93), .ZN(
        \CU_OUTS[EXE][ALU_OP][4] ) );
  AOI22_X1 U115 ( .A1(INSTR_ID[26]), .A2(\CU_OUTS[ID][BRANCH_COND][1] ), .B1(
        \INSTR_ID[27] ), .B2(\CU_OUTS[ID][MUX_IMM_EXT_SEL] ), .ZN(n95) );
  INV_X1 U116 ( .A(n95), .ZN(\CU_OUTS[ID][BRANCH_COND][0] ) );
endmodule


module SNPS_CLOCK_GATE_HIGH_reg_N32_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18782, net18784, net18786, net18787, net18790, net18793;
  assign net18782 = EN;
  assign net18784 = CLK;
  assign ENCLK = net18786;
  assign net18793 = TE;

  DLL_X1 latch ( .D(net18787), .GN(net18784), .Q(net18790) );
  AND2_X1 main_gate ( .A1(net18790), .A2(net18784), .ZN(net18786) );
  OR2_X1 test_or ( .A1(net18782), .A2(net18793), .ZN(net18787) );
endmodule


module reg_N32_0 ( D, EN, CLK, RST, \Q[31] , \Q[30] , \Q[29] , \Q[28] , 
        \Q[27] , \Q[26] , \Q[25] , \Q[24] , \Q[23] , \Q[22] , \Q[21] , \Q[20] , 
        \Q[19] , \Q[18] , \Q[17] , \Q[16] , \Q[15] , \Q[14] , \Q[13] , \Q[12] , 
        \Q[11] , \Q[10] , \Q[9] , \Q[8] , \Q[7] , \Q[6] , \Q[5] , \Q[1] , 
        \Q[0] , \Q[3]_BAR , \Q[2] , \Q[4]_BAR  );
  input [31:0] D;
  input EN, CLK, RST;
  output \Q[31] , \Q[30] , \Q[29] , \Q[28] , \Q[27] , \Q[26] , \Q[25] ,
         \Q[24] , \Q[23] , \Q[22] , \Q[21] , \Q[20] , \Q[19] , \Q[18] ,
         \Q[17] , \Q[16] , \Q[15] , \Q[14] , \Q[13] , \Q[12] , \Q[11] ,
         \Q[10] , \Q[9] , \Q[8] , \Q[7] , \Q[6] , \Q[5] , \Q[1] , \Q[0] ,
         \Q[3]_BAR , \Q[2] , \Q[4]_BAR ;
  wire   net18798, n2;
  wire   [31:0] Q;

  SNPS_CLOCK_GATE_HIGH_reg_N32_0 clk_gate_Q_reg ( .CLK(CLK), .EN(EN), .ENCLK(
        net18798), .TE(1'b0) );
  DFFR_X1 \Q_reg[1]  ( .D(D[1]), .CK(net18798), .RN(RST), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(D[0]), .CK(net18798), .RN(RST), .Q(Q[0]) );
  DFFR_X1 \Q_reg[29]  ( .D(D[29]), .CK(net18798), .RN(RST), .Q(Q[29]) );
  DFFR_X1 \Q_reg[27]  ( .D(D[27]), .CK(net18798), .RN(RST), .Q(Q[27]) );
  DFFR_X1 \Q_reg[31]  ( .D(D[31]), .CK(net18798), .RN(RST), .Q(Q[31]) );
  DFFR_X1 \Q_reg[3]  ( .D(D[3]), .CK(net18798), .RN(RST), .QN(\Q[3]_BAR ) );
  DFFR_X1 \Q_reg[9]  ( .D(D[9]), .CK(net18798), .RN(RST), .Q(Q[9]) );
  DFFR_X1 \Q_reg[8]  ( .D(D[8]), .CK(net18798), .RN(RST), .Q(Q[8]) );
  DFFR_X1 \Q_reg[6]  ( .D(D[6]), .CK(net18798), .RN(RST), .Q(Q[6]) );
  DFFR_X1 \Q_reg[4]  ( .D(D[4]), .CK(net18798), .RN(RST), .QN(\Q[4]_BAR ) );
  DFFR_X1 \Q_reg[7]  ( .D(D[7]), .CK(net18798), .RN(RST), .Q(Q[7]) );
  DFFR_X1 \Q_reg[5]  ( .D(D[5]), .CK(net18798), .RN(RST), .Q(Q[5]) );
  DFFR_X1 \Q_reg[28]  ( .D(D[28]), .CK(net18798), .RN(RST), .Q(Q[28]) );
  DFFR_X1 \Q_reg[26]  ( .D(D[26]), .CK(net18798), .RN(RST), .Q(Q[26]) );
  DFFR_X1 \Q_reg[30]  ( .D(D[30]), .CK(net18798), .RN(RST), .Q(Q[30]) );
  DFFR_X1 \Q_reg[24]  ( .D(D[24]), .CK(net18798), .RN(RST), .Q(Q[24]) );
  DFFR_X1 \Q_reg[13]  ( .D(D[13]), .CK(net18798), .RN(RST), .Q(Q[13]) );
  DFFR_X1 \Q_reg[11]  ( .D(D[11]), .CK(net18798), .RN(RST), .Q(Q[11]) );
  DFFR_X1 \Q_reg[12]  ( .D(D[12]), .CK(net18798), .RN(RST), .Q(Q[12]) );
  DFFR_X1 \Q_reg[10]  ( .D(D[10]), .CK(net18798), .RN(RST), .Q(Q[10]) );
  DFFR_X1 \Q_reg[17]  ( .D(D[17]), .CK(net18798), .RN(RST), .Q(Q[17]) );
  DFFR_X1 \Q_reg[16]  ( .D(D[16]), .CK(net18798), .RN(RST), .Q(Q[16]) );
  DFFR_X1 \Q_reg[15]  ( .D(D[15]), .CK(net18798), .RN(RST), .Q(Q[15]) );
  DFFR_X1 \Q_reg[14]  ( .D(D[14]), .CK(net18798), .RN(RST), .Q(Q[14]) );
  DFFR_X1 \Q_reg[20]  ( .D(D[20]), .CK(net18798), .RN(RST), .Q(Q[20]) );
  DFFR_X1 \Q_reg[19]  ( .D(D[19]), .CK(net18798), .RN(RST), .Q(Q[19]) );
  DFFR_X1 \Q_reg[18]  ( .D(D[18]), .CK(net18798), .RN(RST), .Q(Q[18]) );
  DFFR_X1 \Q_reg[23]  ( .D(D[23]), .CK(net18798), .RN(RST), .Q(Q[23]) );
  DFFR_X1 \Q_reg[22]  ( .D(D[22]), .CK(net18798), .RN(RST), .Q(Q[22]) );
  DFFR_X1 \Q_reg[21]  ( .D(D[21]), .CK(net18798), .RN(RST), .Q(Q[21]) );
  DFFRS_X1 \Q_reg[25]  ( .D(D[25]), .CK(net18798), .RN(RST), .SN(1'b1), .Q(
        Q[25]) );
  DFFS_X1 \Q_reg[2]  ( .D(n2), .CK(net18798), .SN(RST), .QN(Q[2]) );
  INV_X1 U3 ( .A(D[2]), .ZN(n2) );
endmodule


module FA_0 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   A;
  assign S = A;

endmodule


module FA_2079 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   A;
  assign S = A;

endmodule


module FA_2078 ( B, Ci, Co, A, S_BAR );
  input B, Ci, A;
  output Co, S_BAR;
  wire   A;
  assign Co = A;
  assign S_BAR = A;

endmodule


module FA_2077 ( B, Ci, S, Co, A_BAR );
  input B, Ci, A_BAR;
  output S, Co;
  wire   A, n1;
  assign A = A_BAR;

  INV_X1 U1 ( .A(Ci), .ZN(n1) );
  NOR2_X1 U2 ( .A1(A), .A2(n1), .ZN(Co) );
  AOI21_X1 U3 ( .B1(A), .B2(n1), .A(Co), .ZN(S) );
endmodule


module FA_2076 ( B, Ci, S, Co, A_BAR );
  input B, Ci, A_BAR;
  output S, Co;
  wire   A, n1;
  assign A = A_BAR;

  NOR2_X1 U1 ( .A1(A), .A2(n1), .ZN(Co) );
  INV_X1 U2 ( .A(Ci), .ZN(n1) );
  AOI21_X1 U3 ( .B1(A), .B2(n1), .A(Co), .ZN(S) );
endmodule


module FA_2075 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(Ci), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(Ci), .B(A), .Z(S) );
endmodule


module FA_2074 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(Ci), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(Ci), .B(A), .Z(S) );
endmodule


module FA_2073 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(Ci), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(Ci), .B(A), .Z(S) );
endmodule


module FA_2072 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(Ci), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(Ci), .B(A), .Z(S) );
endmodule


module FA_2071 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(Ci), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(Ci), .B(A), .Z(S) );
endmodule


module FA_2070 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(Ci), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(Ci), .B(A), .Z(S) );
endmodule


module FA_2069 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(Ci), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(Ci), .B(A), .Z(S) );
endmodule


module FA_2068 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(Ci), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(Ci), .B(A), .Z(S) );
endmodule


module FA_2067 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(Ci), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(Ci), .B(A), .Z(S) );
endmodule


module FA_2066 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(Ci), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(Ci), .B(A), .Z(S) );
endmodule


module FA_2065 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(Ci), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(Ci), .B(A), .Z(S) );
endmodule


module FA_2064 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(Ci), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(Ci), .B(A), .Z(S) );
endmodule


module FA_2063 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(Ci), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(Ci), .B(A), .Z(S) );
endmodule


module FA_2062 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(Ci), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(Ci), .B(A), .Z(S) );
endmodule


module FA_2061 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(Ci), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(Ci), .B(A), .Z(S) );
endmodule


module FA_2060 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(Ci), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(Ci), .B(A), .Z(S) );
endmodule


module FA_2059 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(Ci), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(Ci), .B(A), .Z(S) );
endmodule


module FA_2058 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(Ci), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(Ci), .B(A), .Z(S) );
endmodule


module FA_2057 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(Ci), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(Ci), .B(A), .Z(S) );
endmodule


module FA_2056 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(Ci), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(Ci), .B(A), .Z(S) );
endmodule


module FA_2055 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(Ci), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(Ci), .B(A), .Z(S) );
endmodule


module FA_2054 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(Ci), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(Ci), .B(A), .Z(S) );
endmodule


module FA_2053 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(Ci), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(Ci), .B(A), .Z(S) );
endmodule


module FA_2052 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(Ci), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(Ci), .B(A), .Z(S) );
endmodule


module FA_2051 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(Ci), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(Ci), .B(A), .Z(S) );
endmodule


module FA_2050 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(Ci), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(Ci), .B(A), .Z(S) );
endmodule


module FA_2049 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XOR2_X1 U1 ( .A(Ci), .B(A), .Z(S) );
endmodule


module RCA_N32 ( B, Ci, Co, \A[31] , \A[30] , \A[29] , \A[28] , \A[27] , 
        \A[26] , \A[25] , \A[24] , \A[23] , \A[22] , \A[21] , \A[20] , \A[19] , 
        \A[18] , \A[17] , \A[16] , \A[15] , \A[14] , \A[13] , \A[12] , \A[11] , 
        \A[10] , \A[9] , \A[8] , \A[7] , \A[6] , \A[5] , \A[1] , \A[0] , 
        \A[3]_BAR , \A[2] , \S[31] , \S[30] , \S[29] , \S[28] , \S[27] , 
        \S[26] , \S[25] , \S[24] , \S[23] , \S[22] , \S[21] , \S[20] , \S[19] , 
        \S[18] , \S[17] , \S[16] , \S[15] , \S[14] , \S[13] , \S[12] , \S[11] , 
        \S[10] , \S[9] , \S[8] , \S[7] , \S[6] , \S[5] , \S[4] , \S[3] , 
        \S[2]_BAR , \S[1] , \S[0] , \A[4]_BAR  );
  input [31:0] B;
  input Ci, \A[31] , \A[30] , \A[29] , \A[28] , \A[27] , \A[26] , \A[25] ,
         \A[24] , \A[23] , \A[22] , \A[21] , \A[20] , \A[19] , \A[18] ,
         \A[17] , \A[16] , \A[15] , \A[14] , \A[13] , \A[12] , \A[11] ,
         \A[10] , \A[9] , \A[8] , \A[7] , \A[6] , \A[5] , \A[1] , \A[0] ,
         \A[3]_BAR , \A[2] , \A[4]_BAR ;
  output Co, \S[31] , \S[30] , \S[29] , \S[28] , \S[27] , \S[26] , \S[25] ,
         \S[24] , \S[23] , \S[22] , \S[21] , \S[20] , \S[19] , \S[18] ,
         \S[17] , \S[16] , \S[15] , \S[14] , \S[13] , \S[12] , \S[11] ,
         \S[10] , \S[9] , \S[8] , \S[7] , \S[6] , \S[5] , \S[4] , \S[3] ,
         \S[2]_BAR , \S[1] , \S[0] ;

  wire   [31:0] A;
  wire   [31:0] S;
  wire   [31:1] CTMP;
  assign A[4] = \A[4]_BAR ;
  assign A[3] = \A[3]_BAR ;
  assign \S[2]_BAR  = S[2];

  FA_0 FULLADDER_1 ( .A(A[0]), .B(1'b0), .Ci(1'b0), .S(S[0]) );
  FA_2079 FULLADDER_2 ( .A(A[1]), .B(1'b0), .Ci(1'b0), .S(S[1]) );
  FA_2078 FULLADDER_3 ( .B(1'b1), .Ci(1'b0), .Co(CTMP[3]), .A(A[2]), .S_BAR(
        S[2]) );
  FA_2077 FULLADDER_4 ( .B(1'b0), .Ci(CTMP[3]), .S(S[3]), .Co(CTMP[4]), 
        .A_BAR(A[3]) );
  FA_2076 FULLADDER_5 ( .B(1'b0), .Ci(CTMP[4]), .S(S[4]), .Co(CTMP[5]), 
        .A_BAR(A[4]) );
  FA_2075 FULLADDER_6 ( .A(A[5]), .B(1'b0), .Ci(CTMP[5]), .S(S[5]), .Co(
        CTMP[6]) );
  FA_2074 FULLADDER_7 ( .A(A[6]), .B(1'b0), .Ci(CTMP[6]), .S(S[6]), .Co(
        CTMP[7]) );
  FA_2073 FULLADDER_8 ( .A(A[7]), .B(1'b0), .Ci(CTMP[7]), .S(S[7]), .Co(
        CTMP[8]) );
  FA_2072 FULLADDER_9 ( .A(A[8]), .B(1'b0), .Ci(CTMP[8]), .S(S[8]), .Co(
        CTMP[9]) );
  FA_2071 FULLADDER_10 ( .A(A[9]), .B(1'b0), .Ci(CTMP[9]), .S(S[9]), .Co(
        CTMP[10]) );
  FA_2070 FULLADDER_11 ( .A(A[10]), .B(1'b0), .Ci(CTMP[10]), .S(S[10]), .Co(
        CTMP[11]) );
  FA_2069 FULLADDER_12 ( .A(A[11]), .B(1'b0), .Ci(CTMP[11]), .S(S[11]), .Co(
        CTMP[12]) );
  FA_2068 FULLADDER_13 ( .A(A[12]), .B(1'b0), .Ci(CTMP[12]), .S(S[12]), .Co(
        CTMP[13]) );
  FA_2067 FULLADDER_14 ( .A(A[13]), .B(1'b0), .Ci(CTMP[13]), .S(S[13]), .Co(
        CTMP[14]) );
  FA_2066 FULLADDER_15 ( .A(A[14]), .B(1'b0), .Ci(CTMP[14]), .S(S[14]), .Co(
        CTMP[15]) );
  FA_2065 FULLADDER_16 ( .A(A[15]), .B(1'b0), .Ci(CTMP[15]), .S(S[15]), .Co(
        CTMP[16]) );
  FA_2064 FULLADDER_17 ( .A(A[16]), .B(1'b0), .Ci(CTMP[16]), .S(S[16]), .Co(
        CTMP[17]) );
  FA_2063 FULLADDER_18 ( .A(A[17]), .B(1'b0), .Ci(CTMP[17]), .S(S[17]), .Co(
        CTMP[18]) );
  FA_2062 FULLADDER_19 ( .A(A[18]), .B(1'b0), .Ci(CTMP[18]), .S(S[18]), .Co(
        CTMP[19]) );
  FA_2061 FULLADDER_20 ( .A(A[19]), .B(1'b0), .Ci(CTMP[19]), .S(S[19]), .Co(
        CTMP[20]) );
  FA_2060 FULLADDER_21 ( .A(A[20]), .B(1'b0), .Ci(CTMP[20]), .S(S[20]), .Co(
        CTMP[21]) );
  FA_2059 FULLADDER_22 ( .A(A[21]), .B(1'b0), .Ci(CTMP[21]), .S(S[21]), .Co(
        CTMP[22]) );
  FA_2058 FULLADDER_23 ( .A(A[22]), .B(1'b0), .Ci(CTMP[22]), .S(S[22]), .Co(
        CTMP[23]) );
  FA_2057 FULLADDER_24 ( .A(A[23]), .B(1'b0), .Ci(CTMP[23]), .S(S[23]), .Co(
        CTMP[24]) );
  FA_2056 FULLADDER_25 ( .A(A[24]), .B(1'b0), .Ci(CTMP[24]), .S(S[24]), .Co(
        CTMP[25]) );
  FA_2055 FULLADDER_26 ( .A(A[25]), .B(1'b0), .Ci(CTMP[25]), .S(S[25]), .Co(
        CTMP[26]) );
  FA_2054 FULLADDER_27 ( .A(A[26]), .B(1'b0), .Ci(CTMP[26]), .S(S[26]), .Co(
        CTMP[27]) );
  FA_2053 FULLADDER_28 ( .A(A[27]), .B(1'b0), .Ci(CTMP[27]), .S(S[27]), .Co(
        CTMP[28]) );
  FA_2052 FULLADDER_29 ( .A(A[28]), .B(1'b0), .Ci(CTMP[28]), .S(S[28]), .Co(
        CTMP[29]) );
  FA_2051 FULLADDER_30 ( .A(A[29]), .B(1'b0), .Ci(CTMP[29]), .S(S[29]), .Co(
        CTMP[30]) );
  FA_2050 FULLADDER_31 ( .A(A[30]), .B(1'b0), .Ci(CTMP[30]), .S(S[30]), .Co(
        CTMP[31]) );
  FA_2049 FULLADDER_32 ( .A(A[31]), .B(1'b0), .Ci(CTMP[31]), .S(S[31]) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_0 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_98 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_97 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_96 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_95 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_94 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_93 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_92 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_91 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_90 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_89 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_88 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_87 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_86 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_85 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_84 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_83 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_82 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_81 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_80 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_79 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_78 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_77 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_76 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_75 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_74 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_73 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_72 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_71 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_70 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_69 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_68 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_67 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_66 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_65 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_64 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_63 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_62 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_61 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_60 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_59 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_58 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_57 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_56 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_55 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_54 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_53 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_52 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_51 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_50 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_49 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_48 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_47 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_46 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_45 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_44 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_43 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_42 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_41 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_40 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_39 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_38 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_37 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_36 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_35 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_34 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_33 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_32 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_31 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_30 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_29 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_28 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_27 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_26 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_25 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_24 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_23 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_22 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_21 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_20 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_19 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_18 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_17 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_16 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_15 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_14 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_13 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_12 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_11 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_10 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_9 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_8 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_7 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_6 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_5 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_4 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_3 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_2 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_1 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net19011, net19013, net19015, net19016, net19019, net19022;
  assign net19011 = EN;
  assign net19013 = CLK;
  assign ENCLK = net19015;
  assign net19022 = TE;

  DLL_X1 latch ( .D(net19016), .GN(net19013), .Q(net19019) );
  AND2_X1 main_gate ( .A1(net19019), .A2(net19013), .ZN(net19015) );
  OR2_X1 test_or ( .A1(net19011), .A2(net19022), .ZN(net19016) );
endmodule


module BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4 ( clk, rst, 
        instr_fetch, pc_out, actual_addr, ID_EN, IF_EN, \pc_fetch[31] , 
        \pc_fetch[30] , \pc_fetch[29] , \pc_fetch[28] , \pc_fetch[27] , 
        \pc_fetch[26] , \pc_fetch[25] , \pc_fetch[24] , \pc_fetch[23] , 
        \pc_fetch[22] , \pc_fetch[21] , \pc_fetch[20] , \pc_fetch[19] , 
        \pc_fetch[18] , \pc_fetch[17] , \pc_fetch[16] , \pc_fetch[15] , 
        \pc_fetch[14] , \pc_fetch[13] , \pc_fetch[12] , \pc_fetch[11] , 
        \pc_fetch[10] , \pc_fetch[9] , \pc_fetch[8] , \pc_fetch[7] , 
        \pc_fetch[6] , \pc_fetch[5] , \pc_fetch[1] , \pc_fetch[0] , 
        \pc_fetch[3]_BAR , misprediction_BAR, \pc_fetch[2] , \pc_in[31] , 
        \pc_in[30] , \pc_in[29] , \pc_in[28] , \pc_in[27] , \pc_in[26] , 
        \pc_in[25] , \pc_in[24] , \pc_in[23] , \pc_in[22] , \pc_in[21] , 
        \pc_in[20] , \pc_in[19] , \pc_in[18] , \pc_in[17] , \pc_in[16] , 
        \pc_in[15] , \pc_in[14] , \pc_in[13] , \pc_in[12] , \pc_in[11] , 
        \pc_in[10] , \pc_in[9] , \pc_in[8] , \pc_in[7] , \pc_in[6] , 
        \pc_in[5] , \pc_in[4] , \pc_in[3] , \pc_in[2]_BAR , \pc_in[1] , 
        \pc_in[0] , \pc_fetch[4]_BAR  );
  input [31:0] instr_fetch;
  output [31:0] pc_out;
  input [31:0] actual_addr;
  input clk, rst, ID_EN, IF_EN, \pc_fetch[31] , \pc_fetch[30] , \pc_fetch[29] ,
         \pc_fetch[28] , \pc_fetch[27] , \pc_fetch[26] , \pc_fetch[25] ,
         \pc_fetch[24] , \pc_fetch[23] , \pc_fetch[22] , \pc_fetch[21] ,
         \pc_fetch[20] , \pc_fetch[19] , \pc_fetch[18] , \pc_fetch[17] ,
         \pc_fetch[16] , \pc_fetch[15] , \pc_fetch[14] , \pc_fetch[13] ,
         \pc_fetch[12] , \pc_fetch[11] , \pc_fetch[10] , \pc_fetch[9] ,
         \pc_fetch[8] , \pc_fetch[7] , \pc_fetch[6] , \pc_fetch[5] ,
         \pc_fetch[1] , \pc_fetch[0] , \pc_fetch[3]_BAR , \pc_fetch[2] ,
         \pc_in[31] , \pc_in[30] , \pc_in[29] , \pc_in[28] , \pc_in[27] ,
         \pc_in[26] , \pc_in[25] , \pc_in[24] , \pc_in[23] , \pc_in[22] ,
         \pc_in[21] , \pc_in[20] , \pc_in[19] , \pc_in[18] , \pc_in[17] ,
         \pc_in[16] , \pc_in[15] , \pc_in[14] , \pc_in[13] , \pc_in[12] ,
         \pc_in[11] , \pc_in[10] , \pc_in[9] , \pc_in[8] , \pc_in[7] ,
         \pc_in[6] , \pc_in[5] , \pc_in[4] , \pc_in[3] , \pc_in[2]_BAR ,
         \pc_in[1] , \pc_in[0] , \pc_fetch[4]_BAR ;
  output misprediction_BAR;
  wire   \hit_index[2] , \hit_index[1] , \hit_index[0] , \cache[0][0][TAG][7] ,
         \cache[0][0][TAG][6] , \cache[0][0][TAG][5] , \cache[0][0][TAG][4] ,
         \cache[0][0][TAG][3] , \cache[0][0][TAG][2] , \cache[0][0][TAG][1] ,
         \cache[0][0][TAG][0] , \cache[0][0][DATA][29] ,
         \cache[0][0][DATA][28] , \cache[0][0][DATA][27] ,
         \cache[0][0][DATA][26] , \cache[0][0][DATA][25] ,
         \cache[0][0][DATA][24] , \cache[0][0][DATA][23] ,
         \cache[0][0][DATA][22] , \cache[0][0][DATA][21] ,
         \cache[0][0][DATA][20] , \cache[0][0][DATA][19] ,
         \cache[0][0][DATA][18] , \cache[0][0][DATA][17] ,
         \cache[0][0][DATA][16] , \cache[0][0][DATA][15] ,
         \cache[0][0][DATA][14] , \cache[0][0][DATA][13] ,
         \cache[0][0][DATA][12] , \cache[0][0][DATA][11] ,
         \cache[0][0][DATA][10] , \cache[0][0][DATA][9] ,
         \cache[0][0][DATA][8] , \cache[0][0][DATA][7] ,
         \cache[0][0][DATA][6] , \cache[0][0][DATA][5] ,
         \cache[0][0][DATA][4] , \cache[0][0][DATA][3] ,
         \cache[0][0][DATA][2] , \cache[0][0][DATA][1] ,
         \cache[0][0][DATA][0] , \cache[0][0][YOUTH][2] ,
         \cache[0][0][YOUTH][1] , \cache[0][0][YOUTH][0] ,
         \cache[0][1][TAG][7] , \cache[0][1][TAG][6] , \cache[0][1][TAG][5] ,
         \cache[0][1][TAG][4] , \cache[0][1][TAG][3] , \cache[0][1][TAG][2] ,
         \cache[0][1][TAG][1] , \cache[0][1][TAG][0] , \cache[0][1][DATA][29] ,
         \cache[0][1][DATA][28] , \cache[0][1][DATA][27] ,
         \cache[0][1][DATA][26] , \cache[0][1][DATA][25] ,
         \cache[0][1][DATA][24] , \cache[0][1][DATA][23] ,
         \cache[0][1][DATA][22] , \cache[0][1][DATA][21] ,
         \cache[0][1][DATA][20] , \cache[0][1][DATA][19] ,
         \cache[0][1][DATA][18] , \cache[0][1][DATA][17] ,
         \cache[0][1][DATA][16] , \cache[0][1][DATA][15] ,
         \cache[0][1][DATA][14] , \cache[0][1][DATA][13] ,
         \cache[0][1][DATA][12] , \cache[0][1][DATA][11] ,
         \cache[0][1][DATA][10] , \cache[0][1][DATA][9] ,
         \cache[0][1][DATA][8] , \cache[0][1][DATA][7] ,
         \cache[0][1][DATA][6] , \cache[0][1][DATA][5] ,
         \cache[0][1][DATA][4] , \cache[0][1][DATA][3] ,
         \cache[0][1][DATA][2] , \cache[0][1][DATA][1] ,
         \cache[0][1][DATA][0] , \cache[0][1][YOUTH][2] ,
         \cache[0][1][YOUTH][1] , \cache[0][1][YOUTH][0] ,
         \cache[0][2][TAG][7] , \cache[0][2][TAG][6] , \cache[0][2][TAG][5] ,
         \cache[0][2][TAG][4] , \cache[0][2][TAG][3] , \cache[0][2][TAG][2] ,
         \cache[0][2][TAG][1] , \cache[0][2][TAG][0] , \cache[0][2][DATA][29] ,
         \cache[0][2][DATA][28] , \cache[0][2][DATA][27] ,
         \cache[0][2][DATA][26] , \cache[0][2][DATA][25] ,
         \cache[0][2][DATA][24] , \cache[0][2][DATA][23] ,
         \cache[0][2][DATA][22] , \cache[0][2][DATA][21] ,
         \cache[0][2][DATA][20] , \cache[0][2][DATA][19] ,
         \cache[0][2][DATA][18] , \cache[0][2][DATA][17] ,
         \cache[0][2][DATA][16] , \cache[0][2][DATA][15] ,
         \cache[0][2][DATA][14] , \cache[0][2][DATA][13] ,
         \cache[0][2][DATA][12] , \cache[0][2][DATA][11] ,
         \cache[0][2][DATA][10] , \cache[0][2][DATA][9] ,
         \cache[0][2][DATA][8] , \cache[0][2][DATA][7] ,
         \cache[0][2][DATA][6] , \cache[0][2][DATA][5] ,
         \cache[0][2][DATA][4] , \cache[0][2][DATA][3] ,
         \cache[0][2][DATA][2] , \cache[0][2][DATA][1] ,
         \cache[0][2][DATA][0] , \cache[0][2][YOUTH][2] ,
         \cache[0][2][YOUTH][1] , \cache[0][2][YOUTH][0] ,
         \cache[0][3][TAG][7] , \cache[0][3][TAG][6] , \cache[0][3][TAG][5] ,
         \cache[0][3][TAG][4] , \cache[0][3][TAG][3] , \cache[0][3][TAG][2] ,
         \cache[0][3][TAG][1] , \cache[0][3][TAG][0] , \cache[0][3][DATA][29] ,
         \cache[0][3][DATA][28] , \cache[0][3][DATA][27] ,
         \cache[0][3][DATA][26] , \cache[0][3][DATA][25] ,
         \cache[0][3][DATA][24] , \cache[0][3][DATA][23] ,
         \cache[0][3][DATA][22] , \cache[0][3][DATA][21] ,
         \cache[0][3][DATA][20] , \cache[0][3][DATA][19] ,
         \cache[0][3][DATA][18] , \cache[0][3][DATA][17] ,
         \cache[0][3][DATA][16] , \cache[0][3][DATA][15] ,
         \cache[0][3][DATA][14] , \cache[0][3][DATA][13] ,
         \cache[0][3][DATA][12] , \cache[0][3][DATA][11] ,
         \cache[0][3][DATA][10] , \cache[0][3][DATA][9] ,
         \cache[0][3][DATA][8] , \cache[0][3][DATA][7] ,
         \cache[0][3][DATA][6] , \cache[0][3][DATA][5] ,
         \cache[0][3][DATA][4] , \cache[0][3][DATA][3] ,
         \cache[0][3][DATA][2] , \cache[0][3][DATA][1] ,
         \cache[0][3][DATA][0] , \cache[0][3][YOUTH][2] ,
         \cache[0][3][YOUTH][1] , \cache[0][3][YOUTH][0] ,
         \cache[1][0][TAG][7] , \cache[1][0][TAG][6] , \cache[1][0][TAG][5] ,
         \cache[1][0][TAG][4] , \cache[1][0][TAG][3] , \cache[1][0][TAG][2] ,
         \cache[1][0][TAG][1] , \cache[1][0][TAG][0] , \cache[1][0][DATA][29] ,
         \cache[1][0][DATA][28] , \cache[1][0][DATA][27] ,
         \cache[1][0][DATA][26] , \cache[1][0][DATA][25] ,
         \cache[1][0][DATA][24] , \cache[1][0][DATA][23] ,
         \cache[1][0][DATA][22] , \cache[1][0][DATA][21] ,
         \cache[1][0][DATA][20] , \cache[1][0][DATA][19] ,
         \cache[1][0][DATA][18] , \cache[1][0][DATA][17] ,
         \cache[1][0][DATA][16] , \cache[1][0][DATA][15] ,
         \cache[1][0][DATA][14] , \cache[1][0][DATA][13] ,
         \cache[1][0][DATA][12] , \cache[1][0][DATA][11] ,
         \cache[1][0][DATA][10] , \cache[1][0][DATA][9] ,
         \cache[1][0][DATA][8] , \cache[1][0][DATA][7] ,
         \cache[1][0][DATA][6] , \cache[1][0][DATA][5] ,
         \cache[1][0][DATA][4] , \cache[1][0][DATA][3] ,
         \cache[1][0][DATA][2] , \cache[1][0][DATA][1] ,
         \cache[1][0][DATA][0] , \cache[1][0][YOUTH][2] ,
         \cache[1][0][YOUTH][1] , \cache[1][0][YOUTH][0] ,
         \cache[1][1][TAG][7] , \cache[1][1][TAG][6] , \cache[1][1][TAG][5] ,
         \cache[1][1][TAG][4] , \cache[1][1][TAG][3] , \cache[1][1][TAG][2] ,
         \cache[1][1][TAG][1] , \cache[1][1][TAG][0] , \cache[1][1][DATA][29] ,
         \cache[1][1][DATA][28] , \cache[1][1][DATA][27] ,
         \cache[1][1][DATA][26] , \cache[1][1][DATA][25] ,
         \cache[1][1][DATA][24] , \cache[1][1][DATA][23] ,
         \cache[1][1][DATA][22] , \cache[1][1][DATA][21] ,
         \cache[1][1][DATA][20] , \cache[1][1][DATA][19] ,
         \cache[1][1][DATA][18] , \cache[1][1][DATA][17] ,
         \cache[1][1][DATA][16] , \cache[1][1][DATA][15] ,
         \cache[1][1][DATA][14] , \cache[1][1][DATA][13] ,
         \cache[1][1][DATA][12] , \cache[1][1][DATA][11] ,
         \cache[1][1][DATA][10] , \cache[1][1][DATA][9] ,
         \cache[1][1][DATA][8] , \cache[1][1][DATA][7] ,
         \cache[1][1][DATA][6] , \cache[1][1][DATA][5] ,
         \cache[1][1][DATA][4] , \cache[1][1][DATA][3] ,
         \cache[1][1][DATA][2] , \cache[1][1][DATA][1] ,
         \cache[1][1][DATA][0] , \cache[1][1][YOUTH][2] ,
         \cache[1][1][YOUTH][1] , \cache[1][1][YOUTH][0] ,
         \cache[1][2][TAG][7] , \cache[1][2][TAG][6] , \cache[1][2][TAG][5] ,
         \cache[1][2][TAG][4] , \cache[1][2][TAG][3] , \cache[1][2][TAG][2] ,
         \cache[1][2][TAG][1] , \cache[1][2][TAG][0] , \cache[1][2][DATA][29] ,
         \cache[1][2][DATA][28] , \cache[1][2][DATA][27] ,
         \cache[1][2][DATA][26] , \cache[1][2][DATA][25] ,
         \cache[1][2][DATA][24] , \cache[1][2][DATA][23] ,
         \cache[1][2][DATA][22] , \cache[1][2][DATA][21] ,
         \cache[1][2][DATA][20] , \cache[1][2][DATA][19] ,
         \cache[1][2][DATA][18] , \cache[1][2][DATA][17] ,
         \cache[1][2][DATA][16] , \cache[1][2][DATA][15] ,
         \cache[1][2][DATA][14] , \cache[1][2][DATA][13] ,
         \cache[1][2][DATA][12] , \cache[1][2][DATA][11] ,
         \cache[1][2][DATA][10] , \cache[1][2][DATA][9] ,
         \cache[1][2][DATA][8] , \cache[1][2][DATA][7] ,
         \cache[1][2][DATA][6] , \cache[1][2][DATA][5] ,
         \cache[1][2][DATA][4] , \cache[1][2][DATA][3] ,
         \cache[1][2][DATA][2] , \cache[1][2][DATA][1] ,
         \cache[1][2][DATA][0] , \cache[1][2][YOUTH][2] ,
         \cache[1][2][YOUTH][1] , \cache[1][2][YOUTH][0] ,
         \cache[1][3][TAG][7] , \cache[1][3][TAG][6] , \cache[1][3][TAG][5] ,
         \cache[1][3][TAG][4] , \cache[1][3][TAG][3] , \cache[1][3][TAG][2] ,
         \cache[1][3][TAG][1] , \cache[1][3][TAG][0] , \cache[1][3][DATA][29] ,
         \cache[1][3][DATA][28] , \cache[1][3][DATA][27] ,
         \cache[1][3][DATA][26] , \cache[1][3][DATA][25] ,
         \cache[1][3][DATA][24] , \cache[1][3][DATA][23] ,
         \cache[1][3][DATA][22] , \cache[1][3][DATA][21] ,
         \cache[1][3][DATA][20] , \cache[1][3][DATA][19] ,
         \cache[1][3][DATA][18] , \cache[1][3][DATA][17] ,
         \cache[1][3][DATA][16] , \cache[1][3][DATA][15] ,
         \cache[1][3][DATA][14] , \cache[1][3][DATA][13] ,
         \cache[1][3][DATA][12] , \cache[1][3][DATA][11] ,
         \cache[1][3][DATA][10] , \cache[1][3][DATA][9] ,
         \cache[1][3][DATA][8] , \cache[1][3][DATA][7] ,
         \cache[1][3][DATA][6] , \cache[1][3][DATA][5] ,
         \cache[1][3][DATA][4] , \cache[1][3][DATA][3] ,
         \cache[1][3][DATA][2] , \cache[1][3][DATA][1] ,
         \cache[1][3][DATA][0] , \cache[1][3][YOUTH][2] ,
         \cache[1][3][YOUTH][1] , \cache[1][3][YOUTH][0] ,
         \cache[2][0][TAG][7] , \cache[2][0][TAG][6] , \cache[2][0][TAG][5] ,
         \cache[2][0][TAG][4] , \cache[2][0][TAG][3] , \cache[2][0][TAG][2] ,
         \cache[2][0][TAG][1] , \cache[2][0][TAG][0] , \cache[2][0][DATA][29] ,
         \cache[2][0][DATA][28] , \cache[2][0][DATA][27] ,
         \cache[2][0][DATA][26] , \cache[2][0][DATA][25] ,
         \cache[2][0][DATA][24] , \cache[2][0][DATA][23] ,
         \cache[2][0][DATA][22] , \cache[2][0][DATA][21] ,
         \cache[2][0][DATA][20] , \cache[2][0][DATA][19] ,
         \cache[2][0][DATA][18] , \cache[2][0][DATA][17] ,
         \cache[2][0][DATA][16] , \cache[2][0][DATA][15] ,
         \cache[2][0][DATA][14] , \cache[2][0][DATA][13] ,
         \cache[2][0][DATA][12] , \cache[2][0][DATA][11] ,
         \cache[2][0][DATA][10] , \cache[2][0][DATA][9] ,
         \cache[2][0][DATA][8] , \cache[2][0][DATA][7] ,
         \cache[2][0][DATA][6] , \cache[2][0][DATA][5] ,
         \cache[2][0][DATA][4] , \cache[2][0][DATA][3] ,
         \cache[2][0][DATA][2] , \cache[2][0][DATA][1] ,
         \cache[2][0][DATA][0] , \cache[2][0][YOUTH][2] ,
         \cache[2][0][YOUTH][1] , \cache[2][0][YOUTH][0] ,
         \cache[2][1][TAG][7] , \cache[2][1][TAG][6] , \cache[2][1][TAG][5] ,
         \cache[2][1][TAG][4] , \cache[2][1][TAG][3] , \cache[2][1][TAG][2] ,
         \cache[2][1][TAG][1] , \cache[2][1][TAG][0] , \cache[2][1][DATA][29] ,
         \cache[2][1][DATA][28] , \cache[2][1][DATA][27] ,
         \cache[2][1][DATA][26] , \cache[2][1][DATA][25] ,
         \cache[2][1][DATA][24] , \cache[2][1][DATA][23] ,
         \cache[2][1][DATA][22] , \cache[2][1][DATA][21] ,
         \cache[2][1][DATA][20] , \cache[2][1][DATA][19] ,
         \cache[2][1][DATA][18] , \cache[2][1][DATA][17] ,
         \cache[2][1][DATA][16] , \cache[2][1][DATA][15] ,
         \cache[2][1][DATA][14] , \cache[2][1][DATA][13] ,
         \cache[2][1][DATA][12] , \cache[2][1][DATA][11] ,
         \cache[2][1][DATA][10] , \cache[2][1][DATA][9] ,
         \cache[2][1][DATA][8] , \cache[2][1][DATA][7] ,
         \cache[2][1][DATA][6] , \cache[2][1][DATA][5] ,
         \cache[2][1][DATA][4] , \cache[2][1][DATA][3] ,
         \cache[2][1][DATA][2] , \cache[2][1][DATA][1] ,
         \cache[2][1][DATA][0] , \cache[2][1][YOUTH][2] ,
         \cache[2][1][YOUTH][1] , \cache[2][1][YOUTH][0] ,
         \cache[2][2][TAG][7] , \cache[2][2][TAG][6] , \cache[2][2][TAG][5] ,
         \cache[2][2][TAG][4] , \cache[2][2][TAG][3] , \cache[2][2][TAG][2] ,
         \cache[2][2][TAG][1] , \cache[2][2][TAG][0] , \cache[2][2][DATA][29] ,
         \cache[2][2][DATA][28] , \cache[2][2][DATA][27] ,
         \cache[2][2][DATA][26] , \cache[2][2][DATA][25] ,
         \cache[2][2][DATA][24] , \cache[2][2][DATA][23] ,
         \cache[2][2][DATA][22] , \cache[2][2][DATA][21] ,
         \cache[2][2][DATA][20] , \cache[2][2][DATA][19] ,
         \cache[2][2][DATA][18] , \cache[2][2][DATA][17] ,
         \cache[2][2][DATA][16] , \cache[2][2][DATA][15] ,
         \cache[2][2][DATA][14] , \cache[2][2][DATA][13] ,
         \cache[2][2][DATA][12] , \cache[2][2][DATA][11] ,
         \cache[2][2][DATA][10] , \cache[2][2][DATA][9] ,
         \cache[2][2][DATA][8] , \cache[2][2][DATA][7] ,
         \cache[2][2][DATA][6] , \cache[2][2][DATA][5] ,
         \cache[2][2][DATA][4] , \cache[2][2][DATA][3] ,
         \cache[2][2][DATA][2] , \cache[2][2][DATA][1] ,
         \cache[2][2][DATA][0] , \cache[2][2][YOUTH][2] ,
         \cache[2][2][YOUTH][1] , \cache[2][2][YOUTH][0] ,
         \cache[2][3][TAG][7] , \cache[2][3][TAG][6] , \cache[2][3][TAG][5] ,
         \cache[2][3][TAG][4] , \cache[2][3][TAG][3] , \cache[2][3][TAG][2] ,
         \cache[2][3][TAG][1] , \cache[2][3][TAG][0] , \cache[2][3][DATA][29] ,
         \cache[2][3][DATA][28] , \cache[2][3][DATA][27] ,
         \cache[2][3][DATA][26] , \cache[2][3][DATA][25] ,
         \cache[2][3][DATA][24] , \cache[2][3][DATA][23] ,
         \cache[2][3][DATA][22] , \cache[2][3][DATA][21] ,
         \cache[2][3][DATA][20] , \cache[2][3][DATA][19] ,
         \cache[2][3][DATA][18] , \cache[2][3][DATA][17] ,
         \cache[2][3][DATA][16] , \cache[2][3][DATA][15] ,
         \cache[2][3][DATA][14] , \cache[2][3][DATA][13] ,
         \cache[2][3][DATA][12] , \cache[2][3][DATA][11] ,
         \cache[2][3][DATA][10] , \cache[2][3][DATA][9] ,
         \cache[2][3][DATA][8] , \cache[2][3][DATA][7] ,
         \cache[2][3][DATA][6] , \cache[2][3][DATA][5] ,
         \cache[2][3][DATA][4] , \cache[2][3][DATA][3] ,
         \cache[2][3][DATA][2] , \cache[2][3][DATA][1] ,
         \cache[2][3][DATA][0] , \cache[2][3][YOUTH][2] ,
         \cache[2][3][YOUTH][1] , \cache[2][3][YOUTH][0] ,
         \cache[3][0][TAG][7] , \cache[3][0][TAG][6] , \cache[3][0][TAG][5] ,
         \cache[3][0][TAG][4] , \cache[3][0][TAG][3] , \cache[3][0][TAG][2] ,
         \cache[3][0][TAG][1] , \cache[3][0][TAG][0] , \cache[3][0][DATA][29] ,
         \cache[3][0][DATA][28] , \cache[3][0][DATA][27] ,
         \cache[3][0][DATA][26] , \cache[3][0][DATA][25] ,
         \cache[3][0][DATA][24] , \cache[3][0][DATA][23] ,
         \cache[3][0][DATA][22] , \cache[3][0][DATA][21] ,
         \cache[3][0][DATA][20] , \cache[3][0][DATA][19] ,
         \cache[3][0][DATA][18] , \cache[3][0][DATA][17] ,
         \cache[3][0][DATA][16] , \cache[3][0][DATA][15] ,
         \cache[3][0][DATA][14] , \cache[3][0][DATA][13] ,
         \cache[3][0][DATA][12] , \cache[3][0][DATA][11] ,
         \cache[3][0][DATA][10] , \cache[3][0][DATA][9] ,
         \cache[3][0][DATA][8] , \cache[3][0][DATA][7] ,
         \cache[3][0][DATA][6] , \cache[3][0][DATA][5] ,
         \cache[3][0][DATA][4] , \cache[3][0][DATA][3] ,
         \cache[3][0][DATA][2] , \cache[3][0][DATA][1] ,
         \cache[3][0][DATA][0] , \cache[3][0][YOUTH][2] ,
         \cache[3][0][YOUTH][1] , \cache[3][0][YOUTH][0] ,
         \cache[3][1][TAG][7] , \cache[3][1][TAG][6] , \cache[3][1][TAG][5] ,
         \cache[3][1][TAG][4] , \cache[3][1][TAG][3] , \cache[3][1][TAG][2] ,
         \cache[3][1][TAG][1] , \cache[3][1][TAG][0] , \cache[3][1][DATA][29] ,
         \cache[3][1][DATA][28] , \cache[3][1][DATA][27] ,
         \cache[3][1][DATA][26] , \cache[3][1][DATA][25] ,
         \cache[3][1][DATA][24] , \cache[3][1][DATA][23] ,
         \cache[3][1][DATA][22] , \cache[3][1][DATA][21] ,
         \cache[3][1][DATA][20] , \cache[3][1][DATA][19] ,
         \cache[3][1][DATA][18] , \cache[3][1][DATA][17] ,
         \cache[3][1][DATA][16] , \cache[3][1][DATA][15] ,
         \cache[3][1][DATA][14] , \cache[3][1][DATA][13] ,
         \cache[3][1][DATA][12] , \cache[3][1][DATA][11] ,
         \cache[3][1][DATA][10] , \cache[3][1][DATA][9] ,
         \cache[3][1][DATA][8] , \cache[3][1][DATA][7] ,
         \cache[3][1][DATA][6] , \cache[3][1][DATA][5] ,
         \cache[3][1][DATA][4] , \cache[3][1][DATA][3] ,
         \cache[3][1][DATA][2] , \cache[3][1][DATA][1] ,
         \cache[3][1][DATA][0] , \cache[3][1][YOUTH][2] ,
         \cache[3][1][YOUTH][1] , \cache[3][1][YOUTH][0] ,
         \cache[3][2][TAG][7] , \cache[3][2][TAG][6] , \cache[3][2][TAG][5] ,
         \cache[3][2][TAG][4] , \cache[3][2][TAG][3] , \cache[3][2][TAG][2] ,
         \cache[3][2][TAG][1] , \cache[3][2][TAG][0] , \cache[3][2][DATA][29] ,
         \cache[3][2][DATA][28] , \cache[3][2][DATA][27] ,
         \cache[3][2][DATA][26] , \cache[3][2][DATA][25] ,
         \cache[3][2][DATA][24] , \cache[3][2][DATA][23] ,
         \cache[3][2][DATA][22] , \cache[3][2][DATA][21] ,
         \cache[3][2][DATA][20] , \cache[3][2][DATA][19] ,
         \cache[3][2][DATA][18] , \cache[3][2][DATA][17] ,
         \cache[3][2][DATA][16] , \cache[3][2][DATA][15] ,
         \cache[3][2][DATA][14] , \cache[3][2][DATA][13] ,
         \cache[3][2][DATA][12] , \cache[3][2][DATA][11] ,
         \cache[3][2][DATA][10] , \cache[3][2][DATA][9] ,
         \cache[3][2][DATA][8] , \cache[3][2][DATA][7] ,
         \cache[3][2][DATA][6] , \cache[3][2][DATA][5] ,
         \cache[3][2][DATA][4] , \cache[3][2][DATA][3] ,
         \cache[3][2][DATA][2] , \cache[3][2][DATA][1] ,
         \cache[3][2][DATA][0] , \cache[3][2][YOUTH][2] ,
         \cache[3][2][YOUTH][1] , \cache[3][2][YOUTH][0] ,
         \cache[3][3][TAG][7] , \cache[3][3][TAG][6] , \cache[3][3][TAG][5] ,
         \cache[3][3][TAG][4] , \cache[3][3][TAG][3] , \cache[3][3][TAG][2] ,
         \cache[3][3][TAG][1] , \cache[3][3][TAG][0] , \cache[3][3][DATA][29] ,
         \cache[3][3][DATA][28] , \cache[3][3][DATA][27] ,
         \cache[3][3][DATA][26] , \cache[3][3][DATA][25] ,
         \cache[3][3][DATA][24] , \cache[3][3][DATA][23] ,
         \cache[3][3][DATA][22] , \cache[3][3][DATA][21] ,
         \cache[3][3][DATA][20] , \cache[3][3][DATA][19] ,
         \cache[3][3][DATA][18] , \cache[3][3][DATA][17] ,
         \cache[3][3][DATA][16] , \cache[3][3][DATA][15] ,
         \cache[3][3][DATA][14] , \cache[3][3][DATA][13] ,
         \cache[3][3][DATA][12] , \cache[3][3][DATA][11] ,
         \cache[3][3][DATA][10] , \cache[3][3][DATA][9] ,
         \cache[3][3][DATA][8] , \cache[3][3][DATA][7] ,
         \cache[3][3][DATA][6] , \cache[3][3][DATA][5] ,
         \cache[3][3][DATA][4] , \cache[3][3][DATA][3] ,
         \cache[3][3][DATA][2] , \cache[3][3][DATA][1] ,
         \cache[3][3][DATA][0] , \cache[3][3][YOUTH][2] ,
         \cache[3][3][YOUTH][1] , \cache[3][3][YOUTH][0] ,
         \cache[4][0][TAG][7] , \cache[4][0][TAG][6] , \cache[4][0][TAG][5] ,
         \cache[4][0][TAG][4] , \cache[4][0][TAG][3] , \cache[4][0][TAG][2] ,
         \cache[4][0][TAG][1] , \cache[4][0][TAG][0] , \cache[4][0][DATA][29] ,
         \cache[4][0][DATA][28] , \cache[4][0][DATA][27] ,
         \cache[4][0][DATA][26] , \cache[4][0][DATA][25] ,
         \cache[4][0][DATA][24] , \cache[4][0][DATA][23] ,
         \cache[4][0][DATA][22] , \cache[4][0][DATA][21] ,
         \cache[4][0][DATA][20] , \cache[4][0][DATA][19] ,
         \cache[4][0][DATA][18] , \cache[4][0][DATA][17] ,
         \cache[4][0][DATA][16] , \cache[4][0][DATA][15] ,
         \cache[4][0][DATA][14] , \cache[4][0][DATA][13] ,
         \cache[4][0][DATA][12] , \cache[4][0][DATA][11] ,
         \cache[4][0][DATA][10] , \cache[4][0][DATA][9] ,
         \cache[4][0][DATA][8] , \cache[4][0][DATA][7] ,
         \cache[4][0][DATA][6] , \cache[4][0][DATA][5] ,
         \cache[4][0][DATA][4] , \cache[4][0][DATA][3] ,
         \cache[4][0][DATA][2] , \cache[4][0][DATA][1] ,
         \cache[4][0][DATA][0] , \cache[4][0][YOUTH][2] ,
         \cache[4][0][YOUTH][1] , \cache[4][0][YOUTH][0] ,
         \cache[4][1][TAG][7] , \cache[4][1][TAG][6] , \cache[4][1][TAG][5] ,
         \cache[4][1][TAG][4] , \cache[4][1][TAG][3] , \cache[4][1][TAG][2] ,
         \cache[4][1][TAG][1] , \cache[4][1][TAG][0] , \cache[4][1][DATA][29] ,
         \cache[4][1][DATA][28] , \cache[4][1][DATA][27] ,
         \cache[4][1][DATA][26] , \cache[4][1][DATA][25] ,
         \cache[4][1][DATA][24] , \cache[4][1][DATA][23] ,
         \cache[4][1][DATA][22] , \cache[4][1][DATA][21] ,
         \cache[4][1][DATA][20] , \cache[4][1][DATA][19] ,
         \cache[4][1][DATA][18] , \cache[4][1][DATA][17] ,
         \cache[4][1][DATA][16] , \cache[4][1][DATA][15] ,
         \cache[4][1][DATA][14] , \cache[4][1][DATA][13] ,
         \cache[4][1][DATA][12] , \cache[4][1][DATA][11] ,
         \cache[4][1][DATA][10] , \cache[4][1][DATA][9] ,
         \cache[4][1][DATA][8] , \cache[4][1][DATA][7] ,
         \cache[4][1][DATA][6] , \cache[4][1][DATA][5] ,
         \cache[4][1][DATA][4] , \cache[4][1][DATA][3] ,
         \cache[4][1][DATA][2] , \cache[4][1][DATA][1] ,
         \cache[4][1][DATA][0] , \cache[4][1][YOUTH][2] ,
         \cache[4][1][YOUTH][1] , \cache[4][1][YOUTH][0] ,
         \cache[4][2][TAG][7] , \cache[4][2][TAG][6] , \cache[4][2][TAG][5] ,
         \cache[4][2][TAG][4] , \cache[4][2][TAG][3] , \cache[4][2][TAG][2] ,
         \cache[4][2][TAG][1] , \cache[4][2][TAG][0] , \cache[4][2][DATA][29] ,
         \cache[4][2][DATA][28] , \cache[4][2][DATA][27] ,
         \cache[4][2][DATA][26] , \cache[4][2][DATA][25] ,
         \cache[4][2][DATA][24] , \cache[4][2][DATA][23] ,
         \cache[4][2][DATA][22] , \cache[4][2][DATA][21] ,
         \cache[4][2][DATA][20] , \cache[4][2][DATA][19] ,
         \cache[4][2][DATA][18] , \cache[4][2][DATA][17] ,
         \cache[4][2][DATA][16] , \cache[4][2][DATA][15] ,
         \cache[4][2][DATA][14] , \cache[4][2][DATA][13] ,
         \cache[4][2][DATA][12] , \cache[4][2][DATA][11] ,
         \cache[4][2][DATA][10] , \cache[4][2][DATA][9] ,
         \cache[4][2][DATA][8] , \cache[4][2][DATA][7] ,
         \cache[4][2][DATA][6] , \cache[4][2][DATA][5] ,
         \cache[4][2][DATA][4] , \cache[4][2][DATA][3] ,
         \cache[4][2][DATA][2] , \cache[4][2][DATA][1] ,
         \cache[4][2][DATA][0] , \cache[4][2][YOUTH][2] ,
         \cache[4][2][YOUTH][1] , \cache[4][2][YOUTH][0] ,
         \cache[4][3][TAG][7] , \cache[4][3][TAG][6] , \cache[4][3][TAG][5] ,
         \cache[4][3][TAG][4] , \cache[4][3][TAG][3] , \cache[4][3][TAG][2] ,
         \cache[4][3][TAG][1] , \cache[4][3][TAG][0] , \cache[4][3][DATA][29] ,
         \cache[4][3][DATA][28] , \cache[4][3][DATA][27] ,
         \cache[4][3][DATA][26] , \cache[4][3][DATA][25] ,
         \cache[4][3][DATA][24] , \cache[4][3][DATA][23] ,
         \cache[4][3][DATA][22] , \cache[4][3][DATA][21] ,
         \cache[4][3][DATA][20] , \cache[4][3][DATA][19] ,
         \cache[4][3][DATA][18] , \cache[4][3][DATA][17] ,
         \cache[4][3][DATA][16] , \cache[4][3][DATA][15] ,
         \cache[4][3][DATA][14] , \cache[4][3][DATA][13] ,
         \cache[4][3][DATA][12] , \cache[4][3][DATA][11] ,
         \cache[4][3][DATA][10] , \cache[4][3][DATA][9] ,
         \cache[4][3][DATA][8] , \cache[4][3][DATA][7] ,
         \cache[4][3][DATA][6] , \cache[4][3][DATA][5] ,
         \cache[4][3][DATA][4] , \cache[4][3][DATA][3] ,
         \cache[4][3][DATA][2] , \cache[4][3][DATA][1] ,
         \cache[4][3][DATA][0] , \cache[4][3][YOUTH][2] ,
         \cache[4][3][YOUTH][1] , \cache[4][3][YOUTH][0] ,
         \cache[5][0][TAG][7] , \cache[5][0][TAG][6] , \cache[5][0][TAG][5] ,
         \cache[5][0][TAG][4] , \cache[5][0][TAG][3] , \cache[5][0][TAG][2] ,
         \cache[5][0][TAG][1] , \cache[5][0][TAG][0] , \cache[5][0][DATA][29] ,
         \cache[5][0][DATA][28] , \cache[5][0][DATA][27] ,
         \cache[5][0][DATA][26] , \cache[5][0][DATA][25] ,
         \cache[5][0][DATA][24] , \cache[5][0][DATA][23] ,
         \cache[5][0][DATA][22] , \cache[5][0][DATA][21] ,
         \cache[5][0][DATA][20] , \cache[5][0][DATA][19] ,
         \cache[5][0][DATA][18] , \cache[5][0][DATA][17] ,
         \cache[5][0][DATA][16] , \cache[5][0][DATA][15] ,
         \cache[5][0][DATA][14] , \cache[5][0][DATA][13] ,
         \cache[5][0][DATA][12] , \cache[5][0][DATA][11] ,
         \cache[5][0][DATA][10] , \cache[5][0][DATA][9] ,
         \cache[5][0][DATA][8] , \cache[5][0][DATA][7] ,
         \cache[5][0][DATA][6] , \cache[5][0][DATA][5] ,
         \cache[5][0][DATA][4] , \cache[5][0][DATA][3] ,
         \cache[5][0][DATA][2] , \cache[5][0][DATA][1] ,
         \cache[5][0][DATA][0] , \cache[5][0][YOUTH][2] ,
         \cache[5][0][YOUTH][1] , \cache[5][0][YOUTH][0] ,
         \cache[5][1][TAG][7] , \cache[5][1][TAG][6] , \cache[5][1][TAG][5] ,
         \cache[5][1][TAG][4] , \cache[5][1][TAG][3] , \cache[5][1][TAG][2] ,
         \cache[5][1][TAG][1] , \cache[5][1][TAG][0] , \cache[5][1][DATA][29] ,
         \cache[5][1][DATA][28] , \cache[5][1][DATA][27] ,
         \cache[5][1][DATA][26] , \cache[5][1][DATA][25] ,
         \cache[5][1][DATA][24] , \cache[5][1][DATA][23] ,
         \cache[5][1][DATA][22] , \cache[5][1][DATA][21] ,
         \cache[5][1][DATA][20] , \cache[5][1][DATA][19] ,
         \cache[5][1][DATA][18] , \cache[5][1][DATA][17] ,
         \cache[5][1][DATA][16] , \cache[5][1][DATA][15] ,
         \cache[5][1][DATA][14] , \cache[5][1][DATA][13] ,
         \cache[5][1][DATA][12] , \cache[5][1][DATA][11] ,
         \cache[5][1][DATA][10] , \cache[5][1][DATA][9] ,
         \cache[5][1][DATA][8] , \cache[5][1][DATA][7] ,
         \cache[5][1][DATA][6] , \cache[5][1][DATA][5] ,
         \cache[5][1][DATA][4] , \cache[5][1][DATA][3] ,
         \cache[5][1][DATA][2] , \cache[5][1][DATA][1] ,
         \cache[5][1][DATA][0] , \cache[5][1][YOUTH][2] ,
         \cache[5][1][YOUTH][1] , \cache[5][1][YOUTH][0] ,
         \cache[5][2][TAG][7] , \cache[5][2][TAG][6] , \cache[5][2][TAG][5] ,
         \cache[5][2][TAG][4] , \cache[5][2][TAG][3] , \cache[5][2][TAG][2] ,
         \cache[5][2][TAG][1] , \cache[5][2][TAG][0] , \cache[5][2][DATA][29] ,
         \cache[5][2][DATA][28] , \cache[5][2][DATA][27] ,
         \cache[5][2][DATA][26] , \cache[5][2][DATA][25] ,
         \cache[5][2][DATA][24] , \cache[5][2][DATA][23] ,
         \cache[5][2][DATA][22] , \cache[5][2][DATA][21] ,
         \cache[5][2][DATA][20] , \cache[5][2][DATA][19] ,
         \cache[5][2][DATA][18] , \cache[5][2][DATA][17] ,
         \cache[5][2][DATA][16] , \cache[5][2][DATA][15] ,
         \cache[5][2][DATA][14] , \cache[5][2][DATA][13] ,
         \cache[5][2][DATA][12] , \cache[5][2][DATA][11] ,
         \cache[5][2][DATA][10] , \cache[5][2][DATA][9] ,
         \cache[5][2][DATA][8] , \cache[5][2][DATA][7] ,
         \cache[5][2][DATA][6] , \cache[5][2][DATA][5] ,
         \cache[5][2][DATA][4] , \cache[5][2][DATA][3] ,
         \cache[5][2][DATA][2] , \cache[5][2][DATA][1] ,
         \cache[5][2][DATA][0] , \cache[5][2][YOUTH][2] ,
         \cache[5][2][YOUTH][1] , \cache[5][2][YOUTH][0] ,
         \cache[5][3][TAG][7] , \cache[5][3][TAG][6] , \cache[5][3][TAG][5] ,
         \cache[5][3][TAG][4] , \cache[5][3][TAG][3] , \cache[5][3][TAG][2] ,
         \cache[5][3][TAG][1] , \cache[5][3][TAG][0] , \cache[5][3][DATA][29] ,
         \cache[5][3][DATA][28] , \cache[5][3][DATA][27] ,
         \cache[5][3][DATA][26] , \cache[5][3][DATA][25] ,
         \cache[5][3][DATA][24] , \cache[5][3][DATA][23] ,
         \cache[5][3][DATA][22] , \cache[5][3][DATA][21] ,
         \cache[5][3][DATA][20] , \cache[5][3][DATA][19] ,
         \cache[5][3][DATA][18] , \cache[5][3][DATA][17] ,
         \cache[5][3][DATA][16] , \cache[5][3][DATA][15] ,
         \cache[5][3][DATA][14] , \cache[5][3][DATA][13] ,
         \cache[5][3][DATA][12] , \cache[5][3][DATA][11] ,
         \cache[5][3][DATA][10] , \cache[5][3][DATA][9] ,
         \cache[5][3][DATA][8] , \cache[5][3][DATA][7] ,
         \cache[5][3][DATA][6] , \cache[5][3][DATA][5] ,
         \cache[5][3][DATA][4] , \cache[5][3][DATA][3] ,
         \cache[5][3][DATA][2] , \cache[5][3][DATA][1] ,
         \cache[5][3][DATA][0] , \cache[5][3][YOUTH][2] ,
         \cache[5][3][YOUTH][1] , \cache[5][3][YOUTH][0] ,
         \cache[6][0][TAG][7] , \cache[6][0][TAG][6] , \cache[6][0][TAG][5] ,
         \cache[6][0][TAG][4] , \cache[6][0][TAG][3] , \cache[6][0][TAG][2] ,
         \cache[6][0][TAG][1] , \cache[6][0][TAG][0] , \cache[6][0][DATA][29] ,
         \cache[6][0][DATA][28] , \cache[6][0][DATA][27] ,
         \cache[6][0][DATA][26] , \cache[6][0][DATA][25] ,
         \cache[6][0][DATA][24] , \cache[6][0][DATA][23] ,
         \cache[6][0][DATA][22] , \cache[6][0][DATA][21] ,
         \cache[6][0][DATA][20] , \cache[6][0][DATA][19] ,
         \cache[6][0][DATA][18] , \cache[6][0][DATA][17] ,
         \cache[6][0][DATA][16] , \cache[6][0][DATA][15] ,
         \cache[6][0][DATA][14] , \cache[6][0][DATA][13] ,
         \cache[6][0][DATA][12] , \cache[6][0][DATA][11] ,
         \cache[6][0][DATA][10] , \cache[6][0][DATA][9] ,
         \cache[6][0][DATA][8] , \cache[6][0][DATA][7] ,
         \cache[6][0][DATA][6] , \cache[6][0][DATA][5] ,
         \cache[6][0][DATA][4] , \cache[6][0][DATA][3] ,
         \cache[6][0][DATA][2] , \cache[6][0][DATA][1] ,
         \cache[6][0][DATA][0] , \cache[6][0][YOUTH][2] ,
         \cache[6][0][YOUTH][1] , \cache[6][0][YOUTH][0] ,
         \cache[6][1][TAG][7] , \cache[6][1][TAG][6] , \cache[6][1][TAG][5] ,
         \cache[6][1][TAG][4] , \cache[6][1][TAG][3] , \cache[6][1][TAG][2] ,
         \cache[6][1][TAG][1] , \cache[6][1][TAG][0] , \cache[6][1][DATA][29] ,
         \cache[6][1][DATA][28] , \cache[6][1][DATA][27] ,
         \cache[6][1][DATA][26] , \cache[6][1][DATA][25] ,
         \cache[6][1][DATA][24] , \cache[6][1][DATA][23] ,
         \cache[6][1][DATA][22] , \cache[6][1][DATA][21] ,
         \cache[6][1][DATA][20] , \cache[6][1][DATA][19] ,
         \cache[6][1][DATA][18] , \cache[6][1][DATA][17] ,
         \cache[6][1][DATA][16] , \cache[6][1][DATA][15] ,
         \cache[6][1][DATA][14] , \cache[6][1][DATA][13] ,
         \cache[6][1][DATA][12] , \cache[6][1][DATA][11] ,
         \cache[6][1][DATA][10] , \cache[6][1][DATA][9] ,
         \cache[6][1][DATA][8] , \cache[6][1][DATA][7] ,
         \cache[6][1][DATA][6] , \cache[6][1][DATA][5] ,
         \cache[6][1][DATA][4] , \cache[6][1][DATA][3] ,
         \cache[6][1][DATA][2] , \cache[6][1][DATA][1] ,
         \cache[6][1][DATA][0] , \cache[6][1][YOUTH][2] ,
         \cache[6][1][YOUTH][1] , \cache[6][1][YOUTH][0] ,
         \cache[6][2][TAG][7] , \cache[6][2][TAG][6] , \cache[6][2][TAG][5] ,
         \cache[6][2][TAG][4] , \cache[6][2][TAG][3] , \cache[6][2][TAG][2] ,
         \cache[6][2][TAG][1] , \cache[6][2][TAG][0] , \cache[6][2][DATA][29] ,
         \cache[6][2][DATA][28] , \cache[6][2][DATA][27] ,
         \cache[6][2][DATA][26] , \cache[6][2][DATA][25] ,
         \cache[6][2][DATA][24] , \cache[6][2][DATA][23] ,
         \cache[6][2][DATA][22] , \cache[6][2][DATA][21] ,
         \cache[6][2][DATA][20] , \cache[6][2][DATA][19] ,
         \cache[6][2][DATA][18] , \cache[6][2][DATA][17] ,
         \cache[6][2][DATA][16] , \cache[6][2][DATA][15] ,
         \cache[6][2][DATA][14] , \cache[6][2][DATA][13] ,
         \cache[6][2][DATA][12] , \cache[6][2][DATA][11] ,
         \cache[6][2][DATA][10] , \cache[6][2][DATA][9] ,
         \cache[6][2][DATA][8] , \cache[6][2][DATA][7] ,
         \cache[6][2][DATA][6] , \cache[6][2][DATA][5] ,
         \cache[6][2][DATA][4] , \cache[6][2][DATA][3] ,
         \cache[6][2][DATA][2] , \cache[6][2][DATA][1] ,
         \cache[6][2][DATA][0] , \cache[6][2][YOUTH][2] ,
         \cache[6][2][YOUTH][1] , \cache[6][2][YOUTH][0] ,
         \cache[6][3][TAG][7] , \cache[6][3][TAG][6] , \cache[6][3][TAG][5] ,
         \cache[6][3][TAG][4] , \cache[6][3][TAG][3] , \cache[6][3][TAG][2] ,
         \cache[6][3][TAG][1] , \cache[6][3][TAG][0] , \cache[6][3][DATA][29] ,
         \cache[6][3][DATA][28] , \cache[6][3][DATA][27] ,
         \cache[6][3][DATA][26] , \cache[6][3][DATA][25] ,
         \cache[6][3][DATA][24] , \cache[6][3][DATA][23] ,
         \cache[6][3][DATA][22] , \cache[6][3][DATA][21] ,
         \cache[6][3][DATA][20] , \cache[6][3][DATA][19] ,
         \cache[6][3][DATA][18] , \cache[6][3][DATA][17] ,
         \cache[6][3][DATA][16] , \cache[6][3][DATA][15] ,
         \cache[6][3][DATA][14] , \cache[6][3][DATA][13] ,
         \cache[6][3][DATA][12] , \cache[6][3][DATA][11] ,
         \cache[6][3][DATA][10] , \cache[6][3][DATA][9] ,
         \cache[6][3][DATA][8] , \cache[6][3][DATA][7] ,
         \cache[6][3][DATA][6] , \cache[6][3][DATA][5] ,
         \cache[6][3][DATA][4] , \cache[6][3][DATA][3] ,
         \cache[6][3][DATA][2] , \cache[6][3][DATA][1] ,
         \cache[6][3][DATA][0] , \cache[6][3][YOUTH][2] ,
         \cache[6][3][YOUTH][1] , \cache[6][3][YOUTH][0] ,
         \cache[7][0][TAG][7] , \cache[7][0][TAG][6] , \cache[7][0][TAG][5] ,
         \cache[7][0][TAG][4] , \cache[7][0][TAG][3] , \cache[7][0][TAG][2] ,
         \cache[7][0][TAG][1] , \cache[7][0][TAG][0] , \cache[7][0][DATA][29] ,
         \cache[7][0][DATA][28] , \cache[7][0][DATA][27] ,
         \cache[7][0][DATA][26] , \cache[7][0][DATA][25] ,
         \cache[7][0][DATA][24] , \cache[7][0][DATA][23] ,
         \cache[7][0][DATA][22] , \cache[7][0][DATA][21] ,
         \cache[7][0][DATA][20] , \cache[7][0][DATA][19] ,
         \cache[7][0][DATA][18] , \cache[7][0][DATA][17] ,
         \cache[7][0][DATA][16] , \cache[7][0][DATA][15] ,
         \cache[7][0][DATA][14] , \cache[7][0][DATA][13] ,
         \cache[7][0][DATA][12] , \cache[7][0][DATA][11] ,
         \cache[7][0][DATA][10] , \cache[7][0][DATA][9] ,
         \cache[7][0][DATA][8] , \cache[7][0][DATA][7] ,
         \cache[7][0][DATA][6] , \cache[7][0][DATA][5] ,
         \cache[7][0][DATA][4] , \cache[7][0][DATA][3] ,
         \cache[7][0][DATA][2] , \cache[7][0][DATA][1] ,
         \cache[7][0][DATA][0] , \cache[7][0][YOUTH][2] ,
         \cache[7][0][YOUTH][1] , \cache[7][0][YOUTH][0] ,
         \cache[7][1][TAG][7] , \cache[7][1][TAG][6] , \cache[7][1][TAG][5] ,
         \cache[7][1][TAG][4] , \cache[7][1][TAG][3] , \cache[7][1][TAG][2] ,
         \cache[7][1][TAG][1] , \cache[7][1][TAG][0] , \cache[7][1][DATA][29] ,
         \cache[7][1][DATA][28] , \cache[7][1][DATA][27] ,
         \cache[7][1][DATA][26] , \cache[7][1][DATA][25] ,
         \cache[7][1][DATA][24] , \cache[7][1][DATA][23] ,
         \cache[7][1][DATA][22] , \cache[7][1][DATA][21] ,
         \cache[7][1][DATA][20] , \cache[7][1][DATA][19] ,
         \cache[7][1][DATA][18] , \cache[7][1][DATA][17] ,
         \cache[7][1][DATA][16] , \cache[7][1][DATA][15] ,
         \cache[7][1][DATA][14] , \cache[7][1][DATA][13] ,
         \cache[7][1][DATA][12] , \cache[7][1][DATA][11] ,
         \cache[7][1][DATA][10] , \cache[7][1][DATA][9] ,
         \cache[7][1][DATA][8] , \cache[7][1][DATA][7] ,
         \cache[7][1][DATA][6] , \cache[7][1][DATA][5] ,
         \cache[7][1][DATA][4] , \cache[7][1][DATA][3] ,
         \cache[7][1][DATA][2] , \cache[7][1][DATA][1] ,
         \cache[7][1][DATA][0] , \cache[7][1][YOUTH][2] ,
         \cache[7][1][YOUTH][1] , \cache[7][1][YOUTH][0] ,
         \cache[7][2][TAG][7] , \cache[7][2][TAG][6] , \cache[7][2][TAG][5] ,
         \cache[7][2][TAG][4] , \cache[7][2][TAG][3] , \cache[7][2][TAG][2] ,
         \cache[7][2][TAG][1] , \cache[7][2][TAG][0] , \cache[7][2][DATA][29] ,
         \cache[7][2][DATA][28] , \cache[7][2][DATA][27] ,
         \cache[7][2][DATA][26] , \cache[7][2][DATA][25] ,
         \cache[7][2][DATA][24] , \cache[7][2][DATA][23] ,
         \cache[7][2][DATA][22] , \cache[7][2][DATA][21] ,
         \cache[7][2][DATA][20] , \cache[7][2][DATA][19] ,
         \cache[7][2][DATA][18] , \cache[7][2][DATA][17] ,
         \cache[7][2][DATA][16] , \cache[7][2][DATA][15] ,
         \cache[7][2][DATA][14] , \cache[7][2][DATA][13] ,
         \cache[7][2][DATA][12] , \cache[7][2][DATA][11] ,
         \cache[7][2][DATA][10] , \cache[7][2][DATA][9] ,
         \cache[7][2][DATA][8] , \cache[7][2][DATA][7] ,
         \cache[7][2][DATA][6] , \cache[7][2][DATA][5] ,
         \cache[7][2][DATA][4] , \cache[7][2][DATA][3] ,
         \cache[7][2][DATA][2] , \cache[7][2][DATA][1] ,
         \cache[7][2][DATA][0] , \cache[7][2][YOUTH][2] ,
         \cache[7][2][YOUTH][1] , \cache[7][2][YOUTH][0] ,
         \cache[7][3][TAG][7] , \cache[7][3][TAG][6] , \cache[7][3][TAG][5] ,
         \cache[7][3][TAG][4] , \cache[7][3][TAG][3] , \cache[7][3][TAG][2] ,
         \cache[7][3][TAG][1] , \cache[7][3][TAG][0] , \cache[7][3][DATA][29] ,
         \cache[7][3][DATA][28] , \cache[7][3][DATA][27] ,
         \cache[7][3][DATA][26] , \cache[7][3][DATA][25] ,
         \cache[7][3][DATA][24] , \cache[7][3][DATA][23] ,
         \cache[7][3][DATA][22] , \cache[7][3][DATA][21] ,
         \cache[7][3][DATA][20] , \cache[7][3][DATA][19] ,
         \cache[7][3][DATA][18] , \cache[7][3][DATA][17] ,
         \cache[7][3][DATA][16] , \cache[7][3][DATA][15] ,
         \cache[7][3][DATA][14] , \cache[7][3][DATA][13] ,
         \cache[7][3][DATA][12] , \cache[7][3][DATA][11] ,
         \cache[7][3][DATA][10] , \cache[7][3][DATA][9] ,
         \cache[7][3][DATA][8] , \cache[7][3][DATA][7] ,
         \cache[7][3][DATA][6] , \cache[7][3][DATA][5] ,
         \cache[7][3][DATA][4] , \cache[7][3][DATA][3] ,
         \cache[7][3][DATA][2] , \cache[7][3][DATA][1] ,
         \cache[7][3][DATA][0] , \cache[7][3][YOUTH][2] ,
         \cache[7][3][YOUTH][1] , \cache[7][3][YOUTH][0] , verify,
         \last_set[2] , \last_set[1] , \last_set[0] , \last_hit_index[2] ,
         \last_hit_index[1] , \last_hit_index[0] , N2805, N2806, N2807, N2811,
         N2812, N2813, N2817, N2818, N2819, N2823, N2824, N2825, N2829, N2830,
         N2831, N2835, N2836, N2837, N2841, N2842, N2843, N2847, N2848, N2849,
         N2853, N2854, N2855, N2859, N2860, N2861, N2865, N2866, N2867, N2871,
         N2872, N2873, N2877, N2878, N2879, N2883, N2884, N2885, N2889, N2890,
         N2891, N2895, N2896, N2897, N2901, N2902, N2903, N2907, N2908, N2909,
         N2913, N2914, N2915, N2919, N2920, N2921, N2925, N2926, N2927, N2931,
         N2932, N2933, N2937, N2938, N2939, N2943, N2944, N2945, N2949, N2950,
         N2951, N2955, N2956, N2957, N2961, N2962, N2963, N2967, N2968, N2969,
         N2973, N2974, N2975, N2979, N2980, N2981, N2985, N2986, N2987, N2991,
         N2992, N2993, N3093, N3094, N3095, N3096, N3097, N3098, N3099, N3100,
         N3101, N3102, N3103, N3104, N3105, N3106, N3107, N3108, N3109, N3110,
         N3111, N3112, N3113, N3114, N3115, N3116, N3117, N3118, N3119, N3120,
         N3121, N3122, N3123, N3124, N3125, N3126, N3127, N3128, N3129, N3130,
         N3131, N3132, N3133, N3134, N3135, N3136, N3137, N3138, N3139, N3140,
         N3141, N3142, N3143, N3144, N3145, N3146, N3147, N3148, N3149, N3150,
         N3151, N3152, N3153, N3154, N3155, N3156, N3157, N3158, N3159, N3160,
         N3161, N3162, N3163, N3164, N3165, N3166, N3167, N3168, N3169, N3170,
         N3171, N3172, N3173, N3174, N3175, N3176, N3177, N3178, N3179, N3180,
         N3181, N3182, N3183, N3184, N3185, N3186, N3187, N3188, N3360, N3361,
         net19027, net19033, net19038, net19043, net19048, net19053, net19058,
         net19063, net19068, net19073, net19078, net19083, net19088, net19093,
         net19098, net19103, net19108, net19113, net19118, net19123, net19128,
         net19133, net19138, net19143, net19148, net19153, net19158, net19163,
         net19168, net19173, net19178, net19183, net19188, net19193, net19198,
         net19203, net19208, net19213, net19218, net19223, net19228, net19233,
         net19238, net19243, net19248, net19253, net19258, net19263, net19268,
         net19273, net19278, net19283, net19288, net19293, net19298, net19303,
         net19308, net19313, net19318, net19323, net19328, net19333, net19338,
         net19343, net19348, net19353, net19358, net19363, net19368, net19373,
         net19378, net19383, net19388, net19393, net19398, net19403, net19408,
         net19413, net19418, net19423, net19428, net19433, net19438, net19443,
         net19448, net19453, net19458, net19463, net19468, net19473, net19478,
         net19483, net19488, net19493, net19498, net19503, net19508, net19513,
         net19518, n1, n2, n3, n4, n5, n6, n7, n8, n64, n65, n66, n67, n585,
         n849, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n55, n56, n57, n58, n59, n60, n61, n62, n63, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586;
  wire   [12:2] pc_fetch;
  wire   [31:0] pc_in;
  wire   [31:0] last_prediction;
  assign pc_fetch[4] = \pc_fetch[4]_BAR ;
  assign pc_fetch[3] = \pc_fetch[3]_BAR ;

  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_0 \clk_gate_cache_reg[0][0][TAG]  ( 
        .CLK(clk), .EN(N3188), .ENCLK(net19027), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_98 \clk_gate_cache_reg[0][0][DATA]  ( 
        .CLK(clk), .EN(N3187), .ENCLK(net19033), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_97 \clk_gate_cache_reg[0][0][YOUTH]  ( 
        .CLK(clk), .EN(N3186), .ENCLK(net19038), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_96 \clk_gate_cache_reg[0][1][TAG]  ( 
        .CLK(clk), .EN(N3185), .ENCLK(net19043), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_95 \clk_gate_cache_reg[0][1][DATA]  ( 
        .CLK(clk), .EN(N3184), .ENCLK(net19048), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_94 \clk_gate_cache_reg[0][1][YOUTH]  ( 
        .CLK(clk), .EN(N3183), .ENCLK(net19053), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_93 \clk_gate_cache_reg[0][2][TAG]  ( 
        .CLK(clk), .EN(N3182), .ENCLK(net19058), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_92 \clk_gate_cache_reg[0][2][DATA]  ( 
        .CLK(clk), .EN(N3181), .ENCLK(net19063), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_91 \clk_gate_cache_reg[0][2][YOUTH]  ( 
        .CLK(clk), .EN(N3180), .ENCLK(net19068), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_90 \clk_gate_cache_reg[0][3][TAG]  ( 
        .CLK(clk), .EN(N3179), .ENCLK(net19073), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_89 \clk_gate_cache_reg[0][3][DATA]  ( 
        .CLK(clk), .EN(N3178), .ENCLK(net19078), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_88 \clk_gate_cache_reg[0][3][YOUTH]  ( 
        .CLK(clk), .EN(N3177), .ENCLK(net19083), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_87 \clk_gate_cache_reg[1][0][TAG]  ( 
        .CLK(clk), .EN(N3176), .ENCLK(net19088), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_86 \clk_gate_cache_reg[1][0][DATA]  ( 
        .CLK(clk), .EN(N3175), .ENCLK(net19093), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_85 \clk_gate_cache_reg[1][0][YOUTH]  ( 
        .CLK(clk), .EN(N3174), .ENCLK(net19098), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_84 \clk_gate_cache_reg[1][1][TAG]  ( 
        .CLK(clk), .EN(N3173), .ENCLK(net19103), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_83 \clk_gate_cache_reg[1][1][DATA]  ( 
        .CLK(clk), .EN(N3172), .ENCLK(net19108), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_82 \clk_gate_cache_reg[1][1][YOUTH]  ( 
        .CLK(clk), .EN(N3171), .ENCLK(net19113), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_81 \clk_gate_cache_reg[1][2][TAG]  ( 
        .CLK(clk), .EN(N3170), .ENCLK(net19118), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_80 \clk_gate_cache_reg[1][2][DATA]  ( 
        .CLK(clk), .EN(N3169), .ENCLK(net19123), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_79 \clk_gate_cache_reg[1][2][YOUTH]  ( 
        .CLK(clk), .EN(N3168), .ENCLK(net19128), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_78 \clk_gate_cache_reg[1][3][TAG]  ( 
        .CLK(clk), .EN(N3167), .ENCLK(net19133), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_77 \clk_gate_cache_reg[1][3][DATA]  ( 
        .CLK(clk), .EN(N3166), .ENCLK(net19138), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_76 \clk_gate_cache_reg[1][3][YOUTH]  ( 
        .CLK(clk), .EN(N3165), .ENCLK(net19143), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_75 \clk_gate_cache_reg[2][0][TAG]  ( 
        .CLK(clk), .EN(N3164), .ENCLK(net19148), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_74 \clk_gate_cache_reg[2][0][DATA]  ( 
        .CLK(clk), .EN(N3163), .ENCLK(net19153), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_73 \clk_gate_cache_reg[2][0][YOUTH]  ( 
        .CLK(clk), .EN(N3162), .ENCLK(net19158), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_72 \clk_gate_cache_reg[2][1][TAG]  ( 
        .CLK(clk), .EN(N3161), .ENCLK(net19163), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_71 \clk_gate_cache_reg[2][1][DATA]  ( 
        .CLK(clk), .EN(N3160), .ENCLK(net19168), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_70 \clk_gate_cache_reg[2][1][YOUTH]  ( 
        .CLK(clk), .EN(N3159), .ENCLK(net19173), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_69 \clk_gate_cache_reg[2][2][TAG]  ( 
        .CLK(clk), .EN(N3158), .ENCLK(net19178), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_68 \clk_gate_cache_reg[2][2][DATA]  ( 
        .CLK(clk), .EN(N3157), .ENCLK(net19183), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_67 \clk_gate_cache_reg[2][2][YOUTH]  ( 
        .CLK(clk), .EN(N3156), .ENCLK(net19188), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_66 \clk_gate_cache_reg[2][3][TAG]  ( 
        .CLK(clk), .EN(N3155), .ENCLK(net19193), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_65 \clk_gate_cache_reg[2][3][DATA]  ( 
        .CLK(clk), .EN(N3154), .ENCLK(net19198), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_64 \clk_gate_cache_reg[2][3][YOUTH]  ( 
        .CLK(clk), .EN(N3153), .ENCLK(net19203), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_63 \clk_gate_cache_reg[3][0][TAG]  ( 
        .CLK(clk), .EN(N3152), .ENCLK(net19208), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_62 \clk_gate_cache_reg[3][0][DATA]  ( 
        .CLK(clk), .EN(N3151), .ENCLK(net19213), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_61 \clk_gate_cache_reg[3][0][YOUTH]  ( 
        .CLK(clk), .EN(N3150), .ENCLK(net19218), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_60 \clk_gate_cache_reg[3][1][TAG]  ( 
        .CLK(clk), .EN(N3149), .ENCLK(net19223), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_59 \clk_gate_cache_reg[3][1][DATA]  ( 
        .CLK(clk), .EN(N3148), .ENCLK(net19228), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_58 \clk_gate_cache_reg[3][1][YOUTH]  ( 
        .CLK(clk), .EN(N3147), .ENCLK(net19233), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_57 \clk_gate_cache_reg[3][2][TAG]  ( 
        .CLK(clk), .EN(N3146), .ENCLK(net19238), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_56 \clk_gate_cache_reg[3][2][DATA]  ( 
        .CLK(clk), .EN(N3145), .ENCLK(net19243), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_55 \clk_gate_cache_reg[3][2][YOUTH]  ( 
        .CLK(clk), .EN(N3144), .ENCLK(net19248), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_54 \clk_gate_cache_reg[3][3][TAG]  ( 
        .CLK(clk), .EN(N3143), .ENCLK(net19253), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_53 \clk_gate_cache_reg[3][3][DATA]  ( 
        .CLK(clk), .EN(N3142), .ENCLK(net19258), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_52 \clk_gate_cache_reg[3][3][YOUTH]  ( 
        .CLK(clk), .EN(N3141), .ENCLK(net19263), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_51 \clk_gate_cache_reg[4][0][TAG]  ( 
        .CLK(clk), .EN(N3140), .ENCLK(net19268), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_50 \clk_gate_cache_reg[4][0][DATA]  ( 
        .CLK(clk), .EN(N3139), .ENCLK(net19273), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_49 \clk_gate_cache_reg[4][0][YOUTH]  ( 
        .CLK(clk), .EN(N3138), .ENCLK(net19278), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_48 \clk_gate_cache_reg[4][1][TAG]  ( 
        .CLK(clk), .EN(N3137), .ENCLK(net19283), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_47 \clk_gate_cache_reg[4][1][DATA]  ( 
        .CLK(clk), .EN(N3136), .ENCLK(net19288), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_46 \clk_gate_cache_reg[4][1][YOUTH]  ( 
        .CLK(clk), .EN(N3135), .ENCLK(net19293), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_45 \clk_gate_cache_reg[4][2][TAG]  ( 
        .CLK(clk), .EN(N3134), .ENCLK(net19298), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_44 \clk_gate_cache_reg[4][2][DATA]  ( 
        .CLK(clk), .EN(N3133), .ENCLK(net19303), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_43 \clk_gate_cache_reg[4][2][YOUTH]  ( 
        .CLK(clk), .EN(N3132), .ENCLK(net19308), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_42 \clk_gate_cache_reg[4][3][TAG]  ( 
        .CLK(clk), .EN(N3131), .ENCLK(net19313), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_41 \clk_gate_cache_reg[4][3][DATA]  ( 
        .CLK(clk), .EN(N3130), .ENCLK(net19318), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_40 \clk_gate_cache_reg[4][3][YOUTH]  ( 
        .CLK(clk), .EN(N3129), .ENCLK(net19323), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_39 \clk_gate_cache_reg[5][0][TAG]  ( 
        .CLK(clk), .EN(N3128), .ENCLK(net19328), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_38 \clk_gate_cache_reg[5][0][DATA]  ( 
        .CLK(clk), .EN(N3127), .ENCLK(net19333), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_37 \clk_gate_cache_reg[5][0][YOUTH]  ( 
        .CLK(clk), .EN(N3126), .ENCLK(net19338), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_36 \clk_gate_cache_reg[5][1][TAG]  ( 
        .CLK(clk), .EN(N3125), .ENCLK(net19343), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_35 \clk_gate_cache_reg[5][1][DATA]  ( 
        .CLK(clk), .EN(N3124), .ENCLK(net19348), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_34 \clk_gate_cache_reg[5][1][YOUTH]  ( 
        .CLK(clk), .EN(N3123), .ENCLK(net19353), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_33 \clk_gate_cache_reg[5][2][TAG]  ( 
        .CLK(clk), .EN(N3122), .ENCLK(net19358), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_32 \clk_gate_cache_reg[5][2][DATA]  ( 
        .CLK(clk), .EN(N3121), .ENCLK(net19363), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_31 \clk_gate_cache_reg[5][2][YOUTH]  ( 
        .CLK(clk), .EN(N3120), .ENCLK(net19368), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_30 \clk_gate_cache_reg[5][3][TAG]  ( 
        .CLK(clk), .EN(N3119), .ENCLK(net19373), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_29 \clk_gate_cache_reg[5][3][DATA]  ( 
        .CLK(clk), .EN(N3118), .ENCLK(net19378), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_28 \clk_gate_cache_reg[5][3][YOUTH]  ( 
        .CLK(clk), .EN(N3117), .ENCLK(net19383), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_27 \clk_gate_cache_reg[6][0][TAG]  ( 
        .CLK(clk), .EN(N3116), .ENCLK(net19388), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_26 \clk_gate_cache_reg[6][0][DATA]  ( 
        .CLK(clk), .EN(N3115), .ENCLK(net19393), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_25 \clk_gate_cache_reg[6][0][YOUTH]  ( 
        .CLK(clk), .EN(N3114), .ENCLK(net19398), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_24 \clk_gate_cache_reg[6][1][TAG]  ( 
        .CLK(clk), .EN(N3113), .ENCLK(net19403), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_23 \clk_gate_cache_reg[6][1][DATA]  ( 
        .CLK(clk), .EN(N3112), .ENCLK(net19408), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_22 \clk_gate_cache_reg[6][1][YOUTH]  ( 
        .CLK(clk), .EN(N3111), .ENCLK(net19413), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_21 \clk_gate_cache_reg[6][2][TAG]  ( 
        .CLK(clk), .EN(N3110), .ENCLK(net19418), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_20 \clk_gate_cache_reg[6][2][DATA]  ( 
        .CLK(clk), .EN(N3109), .ENCLK(net19423), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_19 \clk_gate_cache_reg[6][2][YOUTH]  ( 
        .CLK(clk), .EN(N3108), .ENCLK(net19428), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_18 \clk_gate_cache_reg[6][3][TAG]  ( 
        .CLK(clk), .EN(N3107), .ENCLK(net19433), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_17 \clk_gate_cache_reg[6][3][DATA]  ( 
        .CLK(clk), .EN(N3106), .ENCLK(net19438), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_16 \clk_gate_cache_reg[6][3][YOUTH]  ( 
        .CLK(clk), .EN(N3105), .ENCLK(net19443), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_15 \clk_gate_cache_reg[7][0][TAG]  ( 
        .CLK(clk), .EN(N3104), .ENCLK(net19448), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_14 \clk_gate_cache_reg[7][0][DATA]  ( 
        .CLK(clk), .EN(N3103), .ENCLK(net19453), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_13 \clk_gate_cache_reg[7][0][YOUTH]  ( 
        .CLK(clk), .EN(N3102), .ENCLK(net19458), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_12 \clk_gate_cache_reg[7][1][TAG]  ( 
        .CLK(clk), .EN(N3101), .ENCLK(net19463), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_11 \clk_gate_cache_reg[7][1][DATA]  ( 
        .CLK(clk), .EN(N3100), .ENCLK(net19468), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_10 \clk_gate_cache_reg[7][1][YOUTH]  ( 
        .CLK(clk), .EN(N3099), .ENCLK(net19473), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_9 \clk_gate_cache_reg[7][2][TAG]  ( 
        .CLK(clk), .EN(N3098), .ENCLK(net19478), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_8 \clk_gate_cache_reg[7][2][DATA]  ( 
        .CLK(clk), .EN(N3097), .ENCLK(net19483), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_7 \clk_gate_cache_reg[7][2][YOUTH]  ( 
        .CLK(clk), .EN(N3096), .ENCLK(net19488), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_6 \clk_gate_cache_reg[7][3][TAG]  ( 
        .CLK(clk), .EN(N3095), .ENCLK(net19493), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_5 \clk_gate_cache_reg[7][3][DATA]  ( 
        .CLK(clk), .EN(N3094), .ENCLK(net19498), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_4 \clk_gate_cache_reg[7][3][YOUTH]  ( 
        .CLK(clk), .EN(N3093), .ENCLK(net19503), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_3 clk_gate_verify_reg ( 
        .CLK(clk), .EN(N3360), .ENCLK(net19508), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_2 clk_gate_last_prediction_reg ( 
        .CLK(clk), .EN(N3361), .ENCLK(net19513), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4_1 clk_gate_last_prediction_reg_0 ( 
        .CLK(clk), .EN(N3361), .ENCLK(net19518), .TE(1'b0) );
  DFFS_X1 \last_hit_index_reg[0]  ( .D(\hit_index[0] ), .CK(net19518), .SN(rst), .Q(\last_hit_index[0] ), .QN(n109) );
  DFFS_X1 \cache_reg[7][1][YOUTH][0]  ( .D(N2817), .CK(net19473), .SN(rst), 
        .Q(\cache[7][1][YOUTH][0] ) );
  DFFS_X1 \last_set_reg[2]  ( .D(pc_fetch[4]), .CK(net19518), .SN(rst), .Q(
        n106), .QN(\last_set[2] ) );
  DFFS_X1 \cache_reg[7][1][YOUTH][1]  ( .D(N2818), .CK(net19473), .SN(rst), 
        .Q(\cache[7][1][YOUTH][1] ) );
  DFFS_X1 \last_tag_reg[7]  ( .D(n64), .CK(net19518), .SN(rst), .Q(n8) );
  DFFR_X1 \last_tag_reg[6]  ( .D(pc_fetch[11]), .CK(net19518), .RN(rst), .QN(
        n7) );
  DFFS_X1 \last_tag_reg[5]  ( .D(n65), .CK(net19518), .SN(rst), .Q(n6) );
  DFFR_X1 \last_tag_reg[4]  ( .D(pc_fetch[9]), .CK(net19518), .RN(rst), .QN(n5) );
  DFFS_X1 \last_tag_reg[3]  ( .D(n66), .CK(net19518), .SN(rst), .Q(n4) );
  DFFR_X1 \last_tag_reg[2]  ( .D(pc_fetch[7]), .CK(net19518), .RN(rst), .QN(n3) );
  DFFS_X1 \last_tag_reg[1]  ( .D(n67), .CK(net19518), .SN(rst), .Q(n2) );
  DFFR_X1 \last_tag_reg[0]  ( .D(pc_fetch[5]), .CK(net19518), .RN(rst), .QN(n1) );
  DFFS_X1 \cache_reg[6][1][YOUTH][1]  ( .D(N2842), .CK(net19413), .SN(rst), 
        .Q(\cache[6][1][YOUTH][1] ) );
  DFFS_X1 \cache_reg[6][1][YOUTH][0]  ( .D(N2841), .CK(net19413), .SN(rst), 
        .Q(\cache[6][1][YOUTH][0] ) );
  DFFS_X1 \cache_reg[5][1][YOUTH][1]  ( .D(N2866), .CK(net19353), .SN(rst), 
        .Q(\cache[5][1][YOUTH][1] ) );
  DFFS_X1 \cache_reg[5][1][YOUTH][0]  ( .D(N2865), .CK(net19353), .SN(rst), 
        .Q(\cache[5][1][YOUTH][0] ) );
  DFFS_X1 \cache_reg[4][1][YOUTH][1]  ( .D(N2890), .CK(net19293), .SN(rst), 
        .Q(\cache[4][1][YOUTH][1] ) );
  DFFS_X1 \cache_reg[4][1][YOUTH][0]  ( .D(N2889), .CK(net19293), .SN(rst), 
        .Q(\cache[4][1][YOUTH][0] ) );
  DFFS_X1 \cache_reg[3][1][YOUTH][1]  ( .D(N2914), .CK(net19233), .SN(rst), 
        .Q(\cache[3][1][YOUTH][1] ) );
  DFFS_X1 \cache_reg[3][1][YOUTH][0]  ( .D(N2913), .CK(net19233), .SN(rst), 
        .Q(\cache[3][1][YOUTH][0] ) );
  DFFS_X1 \cache_reg[2][1][YOUTH][1]  ( .D(N2938), .CK(net19173), .SN(rst), 
        .Q(\cache[2][1][YOUTH][1] ) );
  DFFS_X1 \cache_reg[2][1][YOUTH][0]  ( .D(N2937), .CK(net19173), .SN(rst), 
        .Q(\cache[2][1][YOUTH][0] ) );
  DFFS_X1 \cache_reg[1][1][YOUTH][1]  ( .D(N2962), .CK(net19113), .SN(rst), 
        .Q(\cache[1][1][YOUTH][1] ) );
  DFFS_X1 \cache_reg[1][1][YOUTH][0]  ( .D(N2961), .CK(net19113), .SN(rst), 
        .Q(\cache[1][1][YOUTH][0] ) );
  DFFS_X1 \cache_reg[0][1][YOUTH][1]  ( .D(N2986), .CK(net19053), .SN(rst), 
        .Q(\cache[0][1][YOUTH][1] ) );
  DFFS_X1 \cache_reg[0][1][YOUTH][0]  ( .D(N2985), .CK(net19053), .SN(rst), 
        .Q(\cache[0][1][YOUTH][0] ) );
  DFFS_X1 \cache_reg[0][3][YOUTH][0]  ( .D(N2973), .CK(net19083), .SN(rst), 
        .Q(\cache[0][3][YOUTH][0] ) );
  DFFS_X1 \last_hit_index_reg[2]  ( .D(\hit_index[2] ), .CK(net19518), .SN(rst), .Q(\last_hit_index[2] ) );
  DFFS_X1 \cache_reg[0][0][TAG][7]  ( .D(n250), .CK(net19027), .SN(rst), .QN(
        \cache[0][0][TAG][7] ) );
  DFFS_X1 \cache_reg[0][0][TAG][6]  ( .D(n251), .CK(net19027), .SN(rst), .QN(
        \cache[0][0][TAG][6] ) );
  DFFS_X1 \cache_reg[0][0][TAG][5]  ( .D(n252), .CK(net19027), .SN(rst), .QN(
        \cache[0][0][TAG][5] ) );
  DFFS_X1 \cache_reg[0][0][TAG][4]  ( .D(n253), .CK(net19027), .SN(rst), .QN(
        \cache[0][0][TAG][4] ) );
  DFFS_X1 \cache_reg[0][0][TAG][3]  ( .D(n254), .CK(net19027), .SN(rst), .QN(
        \cache[0][0][TAG][3] ) );
  DFFS_X1 \cache_reg[0][0][TAG][2]  ( .D(n255), .CK(net19027), .SN(rst), .QN(
        \cache[0][0][TAG][2] ) );
  DFFS_X1 \cache_reg[0][0][TAG][1]  ( .D(n256), .CK(net19027), .SN(rst), .QN(
        \cache[0][0][TAG][1] ) );
  DFFS_X1 \cache_reg[0][0][TAG][0]  ( .D(n257), .CK(net19027), .SN(rst), .QN(
        \cache[0][0][TAG][0] ) );
  DFFS_X1 \cache_reg[1][0][TAG][7]  ( .D(n8), .CK(net19088), .SN(rst), .QN(
        \cache[1][0][TAG][7] ) );
  DFFS_X1 \cache_reg[1][0][TAG][6]  ( .D(n7), .CK(net19088), .SN(rst), .QN(
        \cache[1][0][TAG][6] ) );
  DFFS_X1 \cache_reg[1][0][TAG][5]  ( .D(n6), .CK(net19088), .SN(rst), .QN(
        \cache[1][0][TAG][5] ) );
  DFFS_X1 \cache_reg[1][0][TAG][4]  ( .D(n5), .CK(net19088), .SN(rst), .QN(
        \cache[1][0][TAG][4] ) );
  DFFS_X1 \cache_reg[1][0][TAG][3]  ( .D(n4), .CK(net19088), .SN(rst), .QN(
        \cache[1][0][TAG][3] ) );
  DFFS_X1 \cache_reg[1][0][TAG][2]  ( .D(n3), .CK(net19088), .SN(rst), .QN(
        \cache[1][0][TAG][2] ) );
  DFFS_X1 \cache_reg[1][0][TAG][1]  ( .D(n2), .CK(net19088), .SN(rst), .QN(
        \cache[1][0][TAG][1] ) );
  DFFS_X1 \cache_reg[1][0][TAG][0]  ( .D(n1), .CK(net19088), .SN(rst), .QN(
        \cache[1][0][TAG][0] ) );
  DFFS_X1 \cache_reg[2][0][TAG][7]  ( .D(n8), .CK(net19148), .SN(rst), .QN(
        \cache[2][0][TAG][7] ) );
  DFFS_X1 \cache_reg[2][0][TAG][6]  ( .D(n7), .CK(net19148), .SN(rst), .QN(
        \cache[2][0][TAG][6] ) );
  DFFS_X1 \cache_reg[2][0][TAG][5]  ( .D(n6), .CK(net19148), .SN(rst), .QN(
        \cache[2][0][TAG][5] ) );
  DFFS_X1 \cache_reg[2][0][TAG][4]  ( .D(n5), .CK(net19148), .SN(n41), .QN(
        \cache[2][0][TAG][4] ) );
  DFFS_X1 \cache_reg[2][0][TAG][3]  ( .D(n4), .CK(net19148), .SN(n41), .QN(
        \cache[2][0][TAG][3] ) );
  DFFS_X1 \cache_reg[2][0][TAG][2]  ( .D(n3), .CK(net19148), .SN(n41), .QN(
        \cache[2][0][TAG][2] ) );
  DFFS_X1 \cache_reg[2][0][TAG][1]  ( .D(n2), .CK(net19148), .SN(n41), .QN(
        \cache[2][0][TAG][1] ) );
  DFFS_X1 \cache_reg[2][0][TAG][0]  ( .D(n1), .CK(net19148), .SN(n41), .QN(
        \cache[2][0][TAG][0] ) );
  DFFS_X1 \cache_reg[3][0][TAG][7]  ( .D(n8), .CK(net19208), .SN(n41), .QN(
        \cache[3][0][TAG][7] ) );
  DFFS_X1 \cache_reg[3][0][TAG][6]  ( .D(n7), .CK(net19208), .SN(n41), .QN(
        \cache[3][0][TAG][6] ) );
  DFFS_X1 \cache_reg[3][0][TAG][5]  ( .D(n6), .CK(net19208), .SN(n41), .QN(
        \cache[3][0][TAG][5] ) );
  DFFS_X1 \cache_reg[3][0][TAG][4]  ( .D(n5), .CK(net19208), .SN(n41), .QN(
        \cache[3][0][TAG][4] ) );
  DFFS_X1 \cache_reg[3][0][TAG][3]  ( .D(n4), .CK(net19208), .SN(n41), .QN(
        \cache[3][0][TAG][3] ) );
  DFFS_X1 \cache_reg[3][0][TAG][2]  ( .D(n3), .CK(net19208), .SN(n41), .QN(
        \cache[3][0][TAG][2] ) );
  DFFS_X1 \cache_reg[3][0][TAG][1]  ( .D(n2), .CK(net19208), .SN(n41), .QN(
        \cache[3][0][TAG][1] ) );
  DFFS_X1 \cache_reg[3][0][TAG][0]  ( .D(n1), .CK(net19208), .SN(n41), .QN(
        \cache[3][0][TAG][0] ) );
  DFFS_X1 \cache_reg[4][0][TAG][7]  ( .D(n8), .CK(net19268), .SN(rst), .QN(
        \cache[4][0][TAG][7] ) );
  DFFS_X1 \cache_reg[4][0][TAG][6]  ( .D(n251), .CK(net19268), .SN(rst), .QN(
        \cache[4][0][TAG][6] ) );
  DFFS_X1 \cache_reg[4][0][TAG][5]  ( .D(n6), .CK(net19268), .SN(rst), .QN(
        \cache[4][0][TAG][5] ) );
  DFFS_X1 \cache_reg[4][0][TAG][4]  ( .D(n253), .CK(net19268), .SN(rst), .QN(
        \cache[4][0][TAG][4] ) );
  DFFS_X1 \cache_reg[4][0][TAG][3]  ( .D(n4), .CK(net19268), .SN(rst), .QN(
        \cache[4][0][TAG][3] ) );
  DFFS_X1 \cache_reg[4][0][TAG][2]  ( .D(n255), .CK(net19268), .SN(rst), .QN(
        \cache[4][0][TAG][2] ) );
  DFFS_X1 \cache_reg[4][0][TAG][1]  ( .D(n2), .CK(net19268), .SN(rst), .QN(
        \cache[4][0][TAG][1] ) );
  DFFS_X1 \cache_reg[4][0][TAG][0]  ( .D(n257), .CK(net19268), .SN(rst), .QN(
        \cache[4][0][TAG][0] ) );
  DFFS_X1 \cache_reg[5][0][TAG][7]  ( .D(n8), .CK(net19328), .SN(rst), .QN(
        \cache[5][0][TAG][7] ) );
  DFFS_X1 \cache_reg[5][0][TAG][6]  ( .D(n7), .CK(net19328), .SN(rst), .QN(
        \cache[5][0][TAG][6] ) );
  DFFS_X1 \cache_reg[5][0][TAG][5]  ( .D(n6), .CK(net19328), .SN(rst), .QN(
        \cache[5][0][TAG][5] ) );
  DFFS_X1 \cache_reg[5][0][TAG][4]  ( .D(n5), .CK(net19328), .SN(rst), .QN(
        \cache[5][0][TAG][4] ) );
  DFFS_X1 \cache_reg[5][0][TAG][3]  ( .D(n4), .CK(net19328), .SN(rst), .QN(
        \cache[5][0][TAG][3] ) );
  DFFS_X1 \cache_reg[5][0][TAG][2]  ( .D(n3), .CK(net19328), .SN(rst), .QN(
        \cache[5][0][TAG][2] ) );
  DFFS_X1 \cache_reg[5][0][TAG][1]  ( .D(n2), .CK(net19328), .SN(rst), .QN(
        \cache[5][0][TAG][1] ) );
  DFFS_X1 \cache_reg[5][0][TAG][0]  ( .D(n1), .CK(net19328), .SN(rst), .QN(
        \cache[5][0][TAG][0] ) );
  DFFS_X1 \cache_reg[6][0][TAG][7]  ( .D(n8), .CK(net19388), .SN(rst), .QN(
        \cache[6][0][TAG][7] ) );
  DFFS_X1 \cache_reg[6][0][TAG][6]  ( .D(n7), .CK(net19388), .SN(rst), .QN(
        \cache[6][0][TAG][6] ) );
  DFFS_X1 \cache_reg[6][0][TAG][5]  ( .D(n6), .CK(net19388), .SN(rst), .QN(
        \cache[6][0][TAG][5] ) );
  DFFS_X1 \cache_reg[6][0][TAG][4]  ( .D(n5), .CK(net19388), .SN(rst), .QN(
        \cache[6][0][TAG][4] ) );
  DFFS_X1 \cache_reg[6][0][TAG][3]  ( .D(n4), .CK(net19388), .SN(rst), .QN(
        \cache[6][0][TAG][3] ) );
  DFFS_X1 \cache_reg[6][0][TAG][2]  ( .D(n3), .CK(net19388), .SN(rst), .QN(
        \cache[6][0][TAG][2] ) );
  DFFS_X1 \cache_reg[6][0][TAG][1]  ( .D(n2), .CK(net19388), .SN(rst), .QN(
        \cache[6][0][TAG][1] ) );
  DFFS_X1 \cache_reg[6][0][TAG][0]  ( .D(n1), .CK(net19388), .SN(rst), .QN(
        \cache[6][0][TAG][0] ) );
  DFFS_X1 \cache_reg[7][0][TAG][7]  ( .D(n8), .CK(net19448), .SN(rst), .QN(
        \cache[7][0][TAG][7] ) );
  DFFS_X1 \cache_reg[7][0][TAG][6]  ( .D(n7), .CK(net19448), .SN(rst), .QN(
        \cache[7][0][TAG][6] ) );
  DFFS_X1 \cache_reg[7][0][TAG][5]  ( .D(n6), .CK(net19448), .SN(rst), .QN(
        \cache[7][0][TAG][5] ) );
  DFFS_X1 \cache_reg[7][0][TAG][4]  ( .D(n5), .CK(net19448), .SN(rst), .QN(
        \cache[7][0][TAG][4] ) );
  DFFS_X1 \cache_reg[7][0][TAG][3]  ( .D(n4), .CK(net19448), .SN(rst), .QN(
        \cache[7][0][TAG][3] ) );
  DFFS_X1 \cache_reg[7][0][TAG][2]  ( .D(n3), .CK(net19448), .SN(rst), .QN(
        \cache[7][0][TAG][2] ) );
  DFFS_X1 \cache_reg[7][0][TAG][1]  ( .D(n2), .CK(net19448), .SN(rst), .QN(
        \cache[7][0][TAG][1] ) );
  DFFS_X1 \cache_reg[7][0][TAG][0]  ( .D(n1), .CK(net19448), .SN(rst), .QN(
        \cache[7][0][TAG][0] ) );
  DFFS_X1 \cache_reg[0][1][TAG][7]  ( .D(n8), .CK(net19043), .SN(rst), .QN(
        \cache[0][1][TAG][7] ) );
  DFFS_X1 \cache_reg[0][1][TAG][6]  ( .D(n7), .CK(net19043), .SN(rst), .QN(
        \cache[0][1][TAG][6] ) );
  DFFS_X1 \cache_reg[0][1][TAG][5]  ( .D(n6), .CK(net19043), .SN(rst), .QN(
        \cache[0][1][TAG][5] ) );
  DFFS_X1 \cache_reg[0][1][TAG][4]  ( .D(n5), .CK(net19043), .SN(rst), .QN(
        \cache[0][1][TAG][4] ) );
  DFFS_X1 \cache_reg[0][1][TAG][3]  ( .D(n4), .CK(net19043), .SN(rst), .QN(
        \cache[0][1][TAG][3] ) );
  DFFS_X1 \cache_reg[0][1][TAG][2]  ( .D(n3), .CK(net19043), .SN(rst), .QN(
        \cache[0][1][TAG][2] ) );
  DFFS_X1 \cache_reg[0][1][TAG][1]  ( .D(n2), .CK(net19043), .SN(rst), .QN(
        \cache[0][1][TAG][1] ) );
  DFFS_X1 \cache_reg[0][1][TAG][0]  ( .D(n1), .CK(net19043), .SN(rst), .QN(
        \cache[0][1][TAG][0] ) );
  DFFS_X1 \cache_reg[1][1][TAG][7]  ( .D(n8), .CK(net19103), .SN(rst), .QN(
        \cache[1][1][TAG][7] ) );
  DFFS_X1 \cache_reg[1][1][TAG][6]  ( .D(n7), .CK(net19103), .SN(rst), .QN(
        \cache[1][1][TAG][6] ) );
  DFFS_X1 \cache_reg[1][1][TAG][5]  ( .D(n6), .CK(net19103), .SN(rst), .QN(
        \cache[1][1][TAG][5] ) );
  DFFS_X1 \cache_reg[1][1][TAG][4]  ( .D(n5), .CK(net19103), .SN(rst), .QN(
        \cache[1][1][TAG][4] ) );
  DFFS_X1 \cache_reg[1][1][TAG][3]  ( .D(n4), .CK(net19103), .SN(n41), .QN(
        \cache[1][1][TAG][3] ) );
  DFFS_X1 \cache_reg[1][1][TAG][2]  ( .D(n3), .CK(net19103), .SN(n41), .QN(
        \cache[1][1][TAG][2] ) );
  DFFS_X1 \cache_reg[1][1][TAG][1]  ( .D(n2), .CK(net19103), .SN(rst), .QN(
        \cache[1][1][TAG][1] ) );
  DFFS_X1 \cache_reg[1][1][TAG][0]  ( .D(n1), .CK(net19103), .SN(rst), .QN(
        \cache[1][1][TAG][0] ) );
  DFFS_X1 \cache_reg[2][1][TAG][7]  ( .D(n8), .CK(net19163), .SN(rst), .QN(
        \cache[2][1][TAG][7] ) );
  DFFS_X1 \cache_reg[2][1][TAG][6]  ( .D(n7), .CK(net19163), .SN(rst), .QN(
        \cache[2][1][TAG][6] ) );
  DFFS_X1 \cache_reg[2][1][TAG][5]  ( .D(n6), .CK(net19163), .SN(rst), .QN(
        \cache[2][1][TAG][5] ) );
  DFFS_X1 \cache_reg[2][1][TAG][4]  ( .D(n5), .CK(net19163), .SN(rst), .QN(
        \cache[2][1][TAG][4] ) );
  DFFS_X1 \cache_reg[2][1][TAG][3]  ( .D(n4), .CK(net19163), .SN(rst), .QN(
        \cache[2][1][TAG][3] ) );
  DFFS_X1 \cache_reg[2][1][TAG][2]  ( .D(n3), .CK(net19163), .SN(rst), .QN(
        \cache[2][1][TAG][2] ) );
  DFFS_X1 \cache_reg[2][1][TAG][1]  ( .D(n2), .CK(net19163), .SN(n41), .QN(
        \cache[2][1][TAG][1] ) );
  DFFS_X1 \cache_reg[2][1][TAG][0]  ( .D(n1), .CK(net19163), .SN(rst), .QN(
        \cache[2][1][TAG][0] ) );
  DFFS_X1 \cache_reg[3][1][TAG][7]  ( .D(n8), .CK(net19223), .SN(n41), .QN(
        \cache[3][1][TAG][7] ) );
  DFFS_X1 \cache_reg[3][1][TAG][6]  ( .D(n7), .CK(net19223), .SN(rst), .QN(
        \cache[3][1][TAG][6] ) );
  DFFS_X1 \cache_reg[3][1][TAG][5]  ( .D(n6), .CK(net19223), .SN(rst), .QN(
        \cache[3][1][TAG][5] ) );
  DFFS_X1 \cache_reg[3][1][TAG][4]  ( .D(n5), .CK(net19223), .SN(rst), .QN(
        \cache[3][1][TAG][4] ) );
  DFFS_X1 \cache_reg[3][1][TAG][3]  ( .D(n4), .CK(net19223), .SN(rst), .QN(
        \cache[3][1][TAG][3] ) );
  DFFS_X1 \cache_reg[3][1][TAG][2]  ( .D(n3), .CK(net19223), .SN(rst), .QN(
        \cache[3][1][TAG][2] ) );
  DFFS_X1 \cache_reg[3][1][TAG][1]  ( .D(n2), .CK(net19223), .SN(n41), .QN(
        \cache[3][1][TAG][1] ) );
  DFFS_X1 \cache_reg[3][1][TAG][0]  ( .D(n1), .CK(net19223), .SN(rst), .QN(
        \cache[3][1][TAG][0] ) );
  DFFS_X1 \cache_reg[4][1][TAG][7]  ( .D(n8), .CK(net19283), .SN(n41), .QN(
        \cache[4][1][TAG][7] ) );
  DFFS_X1 \cache_reg[4][1][TAG][6]  ( .D(n7), .CK(net19283), .SN(rst), .QN(
        \cache[4][1][TAG][6] ) );
  DFFS_X1 \cache_reg[4][1][TAG][5]  ( .D(n6), .CK(net19283), .SN(n41), .QN(
        \cache[4][1][TAG][5] ) );
  DFFS_X1 \cache_reg[4][1][TAG][4]  ( .D(n5), .CK(net19283), .SN(rst), .QN(
        \cache[4][1][TAG][4] ) );
  DFFS_X1 \cache_reg[4][1][TAG][3]  ( .D(n4), .CK(net19283), .SN(rst), .QN(
        \cache[4][1][TAG][3] ) );
  DFFS_X1 \cache_reg[4][1][TAG][2]  ( .D(n3), .CK(net19283), .SN(n41), .QN(
        \cache[4][1][TAG][2] ) );
  DFFS_X1 \cache_reg[4][1][TAG][1]  ( .D(n2), .CK(net19283), .SN(rst), .QN(
        \cache[4][1][TAG][1] ) );
  DFFS_X1 \cache_reg[4][1][TAG][0]  ( .D(n1), .CK(net19283), .SN(rst), .QN(
        \cache[4][1][TAG][0] ) );
  DFFS_X1 \cache_reg[5][1][TAG][7]  ( .D(n8), .CK(net19343), .SN(rst), .QN(
        \cache[5][1][TAG][7] ) );
  DFFS_X1 \cache_reg[5][1][TAG][6]  ( .D(n7), .CK(net19343), .SN(rst), .QN(
        \cache[5][1][TAG][6] ) );
  DFFS_X1 \cache_reg[5][1][TAG][5]  ( .D(n6), .CK(net19343), .SN(rst), .QN(
        \cache[5][1][TAG][5] ) );
  DFFS_X1 \cache_reg[5][1][TAG][4]  ( .D(n5), .CK(net19343), .SN(rst), .QN(
        \cache[5][1][TAG][4] ) );
  DFFS_X1 \cache_reg[5][1][TAG][3]  ( .D(n4), .CK(net19343), .SN(rst), .QN(
        \cache[5][1][TAG][3] ) );
  DFFS_X1 \cache_reg[5][1][TAG][2]  ( .D(n3), .CK(net19343), .SN(rst), .QN(
        \cache[5][1][TAG][2] ) );
  DFFS_X1 \cache_reg[5][1][TAG][1]  ( .D(n2), .CK(net19343), .SN(rst), .QN(
        \cache[5][1][TAG][1] ) );
  DFFS_X1 \cache_reg[5][1][TAG][0]  ( .D(n1), .CK(net19343), .SN(n41), .QN(
        \cache[5][1][TAG][0] ) );
  DFFS_X1 \cache_reg[6][1][TAG][7]  ( .D(n8), .CK(net19403), .SN(rst), .QN(
        \cache[6][1][TAG][7] ) );
  DFFS_X1 \cache_reg[6][1][TAG][6]  ( .D(n7), .CK(net19403), .SN(rst), .QN(
        \cache[6][1][TAG][6] ) );
  DFFS_X1 \cache_reg[6][1][TAG][5]  ( .D(n6), .CK(net19403), .SN(rst), .QN(
        \cache[6][1][TAG][5] ) );
  DFFS_X1 \cache_reg[6][1][TAG][4]  ( .D(n5), .CK(net19403), .SN(n41), .QN(
        \cache[6][1][TAG][4] ) );
  DFFS_X1 \cache_reg[6][1][TAG][3]  ( .D(n4), .CK(net19403), .SN(rst), .QN(
        \cache[6][1][TAG][3] ) );
  DFFS_X1 \cache_reg[6][1][TAG][2]  ( .D(n3), .CK(net19403), .SN(rst), .QN(
        \cache[6][1][TAG][2] ) );
  DFFS_X1 \cache_reg[6][1][TAG][1]  ( .D(n2), .CK(net19403), .SN(rst), .QN(
        \cache[6][1][TAG][1] ) );
  DFFS_X1 \cache_reg[6][1][TAG][0]  ( .D(n1), .CK(net19403), .SN(rst), .QN(
        \cache[6][1][TAG][0] ) );
  DFFS_X1 \cache_reg[7][1][TAG][7]  ( .D(n8), .CK(net19463), .SN(rst), .QN(
        \cache[7][1][TAG][7] ) );
  DFFS_X1 \cache_reg[7][1][TAG][6]  ( .D(n7), .CK(net19463), .SN(rst), .QN(
        \cache[7][1][TAG][6] ) );
  DFFS_X1 \cache_reg[7][1][TAG][5]  ( .D(n6), .CK(net19463), .SN(rst), .QN(
        \cache[7][1][TAG][5] ) );
  DFFS_X1 \cache_reg[7][1][TAG][4]  ( .D(n5), .CK(net19463), .SN(rst), .QN(
        \cache[7][1][TAG][4] ) );
  DFFS_X1 \cache_reg[7][1][TAG][3]  ( .D(n4), .CK(net19463), .SN(rst), .QN(
        \cache[7][1][TAG][3] ) );
  DFFS_X1 \cache_reg[7][1][TAG][2]  ( .D(n3), .CK(net19463), .SN(rst), .QN(
        \cache[7][1][TAG][2] ) );
  DFFS_X1 \cache_reg[7][1][TAG][1]  ( .D(n2), .CK(net19463), .SN(rst), .QN(
        \cache[7][1][TAG][1] ) );
  DFFS_X1 \cache_reg[7][1][TAG][0]  ( .D(n1), .CK(net19463), .SN(rst), .QN(
        \cache[7][1][TAG][0] ) );
  DFFS_X1 \cache_reg[0][2][TAG][7]  ( .D(n8), .CK(net19058), .SN(rst), .QN(
        \cache[0][2][TAG][7] ) );
  DFFS_X1 \cache_reg[0][2][TAG][6]  ( .D(n7), .CK(net19058), .SN(rst), .QN(
        \cache[0][2][TAG][6] ) );
  DFFS_X1 \cache_reg[0][2][TAG][5]  ( .D(n6), .CK(net19058), .SN(rst), .QN(
        \cache[0][2][TAG][5] ) );
  DFFS_X1 \cache_reg[0][2][TAG][4]  ( .D(n5), .CK(net19058), .SN(rst), .QN(
        \cache[0][2][TAG][4] ) );
  DFFS_X1 \cache_reg[0][2][TAG][3]  ( .D(n4), .CK(net19058), .SN(rst), .QN(
        \cache[0][2][TAG][3] ) );
  DFFS_X1 \cache_reg[0][2][TAG][2]  ( .D(n3), .CK(net19058), .SN(rst), .QN(
        \cache[0][2][TAG][2] ) );
  DFFS_X1 \cache_reg[0][2][TAG][1]  ( .D(n2), .CK(net19058), .SN(rst), .QN(
        \cache[0][2][TAG][1] ) );
  DFFS_X1 \cache_reg[0][2][TAG][0]  ( .D(n1), .CK(net19058), .SN(rst), .QN(
        \cache[0][2][TAG][0] ) );
  DFFS_X1 \cache_reg[1][2][TAG][7]  ( .D(n8), .CK(net19118), .SN(rst), .QN(
        \cache[1][2][TAG][7] ) );
  DFFS_X1 \cache_reg[1][2][TAG][6]  ( .D(n7), .CK(net19118), .SN(rst), .QN(
        \cache[1][2][TAG][6] ) );
  DFFS_X1 \cache_reg[1][2][TAG][5]  ( .D(n6), .CK(net19118), .SN(rst), .QN(
        \cache[1][2][TAG][5] ) );
  DFFS_X1 \cache_reg[1][2][TAG][4]  ( .D(n5), .CK(net19118), .SN(rst), .QN(
        \cache[1][2][TAG][4] ) );
  DFFS_X1 \cache_reg[1][2][TAG][3]  ( .D(n4), .CK(net19118), .SN(rst), .QN(
        \cache[1][2][TAG][3] ) );
  DFFS_X1 \cache_reg[1][2][TAG][2]  ( .D(n3), .CK(net19118), .SN(rst), .QN(
        \cache[1][2][TAG][2] ) );
  DFFS_X1 \cache_reg[1][2][TAG][1]  ( .D(n2), .CK(net19118), .SN(rst), .QN(
        \cache[1][2][TAG][1] ) );
  DFFS_X1 \cache_reg[1][2][TAG][0]  ( .D(n1), .CK(net19118), .SN(rst), .QN(
        \cache[1][2][TAG][0] ) );
  DFFS_X1 \cache_reg[2][2][TAG][7]  ( .D(n8), .CK(net19178), .SN(rst), .QN(
        \cache[2][2][TAG][7] ) );
  DFFS_X1 \cache_reg[2][2][TAG][6]  ( .D(n7), .CK(net19178), .SN(rst), .QN(
        \cache[2][2][TAG][6] ) );
  DFFS_X1 \cache_reg[2][2][TAG][5]  ( .D(n6), .CK(net19178), .SN(rst), .QN(
        \cache[2][2][TAG][5] ) );
  DFFS_X1 \cache_reg[2][2][TAG][4]  ( .D(n5), .CK(net19178), .SN(rst), .QN(
        \cache[2][2][TAG][4] ) );
  DFFS_X1 \cache_reg[2][2][TAG][3]  ( .D(n4), .CK(net19178), .SN(rst), .QN(
        \cache[2][2][TAG][3] ) );
  DFFS_X1 \cache_reg[2][2][TAG][2]  ( .D(n3), .CK(net19178), .SN(rst), .QN(
        \cache[2][2][TAG][2] ) );
  DFFS_X1 \cache_reg[2][2][TAG][1]  ( .D(n2), .CK(net19178), .SN(rst), .QN(
        \cache[2][2][TAG][1] ) );
  DFFS_X1 \cache_reg[2][2][TAG][0]  ( .D(n1), .CK(net19178), .SN(rst), .QN(
        \cache[2][2][TAG][0] ) );
  DFFS_X1 \cache_reg[3][2][TAG][7]  ( .D(n8), .CK(net19238), .SN(rst), .QN(
        \cache[3][2][TAG][7] ) );
  DFFS_X1 \cache_reg[3][2][TAG][6]  ( .D(n7), .CK(net19238), .SN(rst), .QN(
        \cache[3][2][TAG][6] ) );
  DFFS_X1 \cache_reg[3][2][TAG][5]  ( .D(n6), .CK(net19238), .SN(rst), .QN(
        \cache[3][2][TAG][5] ) );
  DFFS_X1 \cache_reg[3][2][TAG][4]  ( .D(n5), .CK(net19238), .SN(rst), .QN(
        \cache[3][2][TAG][4] ) );
  DFFS_X1 \cache_reg[3][2][TAG][3]  ( .D(n4), .CK(net19238), .SN(rst), .QN(
        \cache[3][2][TAG][3] ) );
  DFFS_X1 \cache_reg[3][2][TAG][2]  ( .D(n3), .CK(net19238), .SN(rst), .QN(
        \cache[3][2][TAG][2] ) );
  DFFS_X1 \cache_reg[3][2][TAG][1]  ( .D(n2), .CK(net19238), .SN(rst), .QN(
        \cache[3][2][TAG][1] ) );
  DFFS_X1 \cache_reg[3][2][TAG][0]  ( .D(n1), .CK(net19238), .SN(rst), .QN(
        \cache[3][2][TAG][0] ) );
  DFFS_X1 \cache_reg[4][2][TAG][7]  ( .D(n8), .CK(net19298), .SN(rst), .QN(
        \cache[4][2][TAG][7] ) );
  DFFS_X1 \cache_reg[4][2][TAG][6]  ( .D(n7), .CK(net19298), .SN(rst), .QN(
        \cache[4][2][TAG][6] ) );
  DFFS_X1 \cache_reg[4][2][TAG][5]  ( .D(n6), .CK(net19298), .SN(rst), .QN(
        \cache[4][2][TAG][5] ) );
  DFFS_X1 \cache_reg[4][2][TAG][4]  ( .D(n5), .CK(net19298), .SN(rst), .QN(
        \cache[4][2][TAG][4] ) );
  DFFS_X1 \cache_reg[4][2][TAG][3]  ( .D(n4), .CK(net19298), .SN(rst), .QN(
        \cache[4][2][TAG][3] ) );
  DFFS_X1 \cache_reg[4][2][TAG][2]  ( .D(n3), .CK(net19298), .SN(rst), .QN(
        \cache[4][2][TAG][2] ) );
  DFFS_X1 \cache_reg[4][2][TAG][1]  ( .D(n2), .CK(net19298), .SN(rst), .QN(
        \cache[4][2][TAG][1] ) );
  DFFS_X1 \cache_reg[4][2][TAG][0]  ( .D(n1), .CK(net19298), .SN(rst), .QN(
        \cache[4][2][TAG][0] ) );
  DFFS_X1 \cache_reg[5][2][TAG][7]  ( .D(n8), .CK(net19358), .SN(rst), .QN(
        \cache[5][2][TAG][7] ) );
  DFFS_X1 \cache_reg[5][2][TAG][6]  ( .D(n7), .CK(net19358), .SN(rst), .QN(
        \cache[5][2][TAG][6] ) );
  DFFS_X1 \cache_reg[5][2][TAG][5]  ( .D(n6), .CK(net19358), .SN(rst), .QN(
        \cache[5][2][TAG][5] ) );
  DFFS_X1 \cache_reg[5][2][TAG][4]  ( .D(n5), .CK(net19358), .SN(rst), .QN(
        \cache[5][2][TAG][4] ) );
  DFFS_X1 \cache_reg[5][2][TAG][3]  ( .D(n4), .CK(net19358), .SN(rst), .QN(
        \cache[5][2][TAG][3] ) );
  DFFS_X1 \cache_reg[5][2][TAG][2]  ( .D(n3), .CK(net19358), .SN(rst), .QN(
        \cache[5][2][TAG][2] ) );
  DFFS_X1 \cache_reg[5][2][TAG][1]  ( .D(n2), .CK(net19358), .SN(rst), .QN(
        \cache[5][2][TAG][1] ) );
  DFFS_X1 \cache_reg[5][2][TAG][0]  ( .D(n1), .CK(net19358), .SN(rst), .QN(
        \cache[5][2][TAG][0] ) );
  DFFS_X1 \cache_reg[6][2][TAG][7]  ( .D(n250), .CK(net19418), .SN(rst), .QN(
        \cache[6][2][TAG][7] ) );
  DFFS_X1 \cache_reg[6][2][TAG][6]  ( .D(n251), .CK(net19418), .SN(rst), .QN(
        \cache[6][2][TAG][6] ) );
  DFFS_X1 \cache_reg[6][2][TAG][5]  ( .D(n252), .CK(net19418), .SN(rst), .QN(
        \cache[6][2][TAG][5] ) );
  DFFS_X1 \cache_reg[6][2][TAG][4]  ( .D(n253), .CK(net19418), .SN(rst), .QN(
        \cache[6][2][TAG][4] ) );
  DFFS_X1 \cache_reg[6][2][TAG][3]  ( .D(n254), .CK(net19418), .SN(rst), .QN(
        \cache[6][2][TAG][3] ) );
  DFFS_X1 \cache_reg[6][2][TAG][2]  ( .D(n255), .CK(net19418), .SN(rst), .QN(
        \cache[6][2][TAG][2] ) );
  DFFS_X1 \cache_reg[6][2][TAG][1]  ( .D(n256), .CK(net19418), .SN(rst), .QN(
        \cache[6][2][TAG][1] ) );
  DFFS_X1 \cache_reg[6][2][TAG][0]  ( .D(n257), .CK(net19418), .SN(rst), .QN(
        \cache[6][2][TAG][0] ) );
  DFFS_X1 \cache_reg[7][2][TAG][7]  ( .D(n250), .CK(net19478), .SN(rst), .QN(
        \cache[7][2][TAG][7] ) );
  DFFS_X1 \cache_reg[7][2][TAG][6]  ( .D(n251), .CK(net19478), .SN(rst), .QN(
        \cache[7][2][TAG][6] ) );
  DFFS_X1 \cache_reg[7][2][TAG][5]  ( .D(n252), .CK(net19478), .SN(rst), .QN(
        \cache[7][2][TAG][5] ) );
  DFFS_X1 \cache_reg[7][2][TAG][4]  ( .D(n253), .CK(net19478), .SN(rst), .QN(
        \cache[7][2][TAG][4] ) );
  DFFS_X1 \cache_reg[7][2][TAG][3]  ( .D(n254), .CK(net19478), .SN(rst), .QN(
        \cache[7][2][TAG][3] ) );
  DFFS_X1 \cache_reg[7][2][TAG][2]  ( .D(n255), .CK(net19478), .SN(rst), .QN(
        \cache[7][2][TAG][2] ) );
  DFFS_X1 \cache_reg[7][2][TAG][1]  ( .D(n256), .CK(net19478), .SN(rst), .QN(
        \cache[7][2][TAG][1] ) );
  DFFS_X1 \cache_reg[7][2][TAG][0]  ( .D(n257), .CK(net19478), .SN(rst), .QN(
        \cache[7][2][TAG][0] ) );
  DFFS_X1 \cache_reg[0][3][TAG][7]  ( .D(n250), .CK(net19073), .SN(rst), .QN(
        \cache[0][3][TAG][7] ) );
  DFFS_X1 \cache_reg[0][3][TAG][6]  ( .D(n251), .CK(net19073), .SN(rst), .QN(
        \cache[0][3][TAG][6] ) );
  DFFS_X1 \cache_reg[0][3][TAG][5]  ( .D(n252), .CK(net19073), .SN(rst), .QN(
        \cache[0][3][TAG][5] ) );
  DFFS_X1 \cache_reg[0][3][TAG][4]  ( .D(n253), .CK(net19073), .SN(rst), .QN(
        \cache[0][3][TAG][4] ) );
  DFFS_X1 \cache_reg[0][3][TAG][3]  ( .D(n254), .CK(net19073), .SN(rst), .QN(
        \cache[0][3][TAG][3] ) );
  DFFS_X1 \cache_reg[0][3][TAG][2]  ( .D(n255), .CK(net19073), .SN(rst), .QN(
        \cache[0][3][TAG][2] ) );
  DFFS_X1 \cache_reg[0][3][TAG][1]  ( .D(n256), .CK(net19073), .SN(rst), .QN(
        \cache[0][3][TAG][1] ) );
  DFFS_X1 \cache_reg[0][3][TAG][0]  ( .D(n257), .CK(net19073), .SN(rst), .QN(
        \cache[0][3][TAG][0] ) );
  DFFS_X1 \cache_reg[1][3][TAG][7]  ( .D(n250), .CK(net19133), .SN(rst), .QN(
        \cache[1][3][TAG][7] ) );
  DFFS_X1 \cache_reg[1][3][TAG][6]  ( .D(n251), .CK(net19133), .SN(rst), .QN(
        \cache[1][3][TAG][6] ) );
  DFFS_X1 \cache_reg[1][3][TAG][5]  ( .D(n252), .CK(net19133), .SN(rst), .QN(
        \cache[1][3][TAG][5] ) );
  DFFS_X1 \cache_reg[1][3][TAG][4]  ( .D(n253), .CK(net19133), .SN(rst), .QN(
        \cache[1][3][TAG][4] ) );
  DFFS_X1 \cache_reg[1][3][TAG][3]  ( .D(n254), .CK(net19133), .SN(rst), .QN(
        \cache[1][3][TAG][3] ) );
  DFFS_X1 \cache_reg[1][3][TAG][2]  ( .D(n255), .CK(net19133), .SN(rst), .QN(
        \cache[1][3][TAG][2] ) );
  DFFS_X1 \cache_reg[1][3][TAG][1]  ( .D(n256), .CK(net19133), .SN(rst), .QN(
        \cache[1][3][TAG][1] ) );
  DFFS_X1 \cache_reg[1][3][TAG][0]  ( .D(n257), .CK(net19133), .SN(rst), .QN(
        \cache[1][3][TAG][0] ) );
  DFFS_X1 \cache_reg[2][3][TAG][7]  ( .D(n250), .CK(net19193), .SN(rst), .QN(
        \cache[2][3][TAG][7] ) );
  DFFS_X1 \cache_reg[2][3][TAG][6]  ( .D(n251), .CK(net19193), .SN(rst), .QN(
        \cache[2][3][TAG][6] ) );
  DFFS_X1 \cache_reg[2][3][TAG][5]  ( .D(n252), .CK(net19193), .SN(rst), .QN(
        \cache[2][3][TAG][5] ) );
  DFFS_X1 \cache_reg[2][3][TAG][4]  ( .D(n253), .CK(net19193), .SN(rst), .QN(
        \cache[2][3][TAG][4] ) );
  DFFS_X1 \cache_reg[2][3][TAG][3]  ( .D(n254), .CK(net19193), .SN(rst), .QN(
        \cache[2][3][TAG][3] ) );
  DFFS_X1 \cache_reg[2][3][TAG][2]  ( .D(n255), .CK(net19193), .SN(rst), .QN(
        \cache[2][3][TAG][2] ) );
  DFFS_X1 \cache_reg[2][3][TAG][1]  ( .D(n256), .CK(net19193), .SN(rst), .QN(
        \cache[2][3][TAG][1] ) );
  DFFS_X1 \cache_reg[2][3][TAG][0]  ( .D(n257), .CK(net19193), .SN(rst), .QN(
        \cache[2][3][TAG][0] ) );
  DFFS_X1 \cache_reg[3][3][TAG][7]  ( .D(n250), .CK(net19253), .SN(rst), .QN(
        \cache[3][3][TAG][7] ) );
  DFFS_X1 \cache_reg[3][3][TAG][6]  ( .D(n251), .CK(net19253), .SN(rst), .QN(
        \cache[3][3][TAG][6] ) );
  DFFS_X1 \cache_reg[3][3][TAG][5]  ( .D(n252), .CK(net19253), .SN(rst), .QN(
        \cache[3][3][TAG][5] ) );
  DFFS_X1 \cache_reg[3][3][TAG][4]  ( .D(n253), .CK(net19253), .SN(rst), .QN(
        \cache[3][3][TAG][4] ) );
  DFFS_X1 \cache_reg[3][3][TAG][3]  ( .D(n254), .CK(net19253), .SN(rst), .QN(
        \cache[3][3][TAG][3] ) );
  DFFS_X1 \cache_reg[3][3][TAG][2]  ( .D(n255), .CK(net19253), .SN(rst), .QN(
        \cache[3][3][TAG][2] ) );
  DFFS_X1 \cache_reg[3][3][TAG][1]  ( .D(n256), .CK(net19253), .SN(rst), .QN(
        \cache[3][3][TAG][1] ) );
  DFFS_X1 \cache_reg[3][3][TAG][0]  ( .D(n257), .CK(net19253), .SN(rst), .QN(
        \cache[3][3][TAG][0] ) );
  DFFS_X1 \cache_reg[4][3][TAG][7]  ( .D(n250), .CK(net19313), .SN(rst), .QN(
        \cache[4][3][TAG][7] ) );
  DFFS_X1 \cache_reg[4][3][TAG][6]  ( .D(n251), .CK(net19313), .SN(rst), .QN(
        \cache[4][3][TAG][6] ) );
  DFFS_X1 \cache_reg[4][3][TAG][5]  ( .D(n252), .CK(net19313), .SN(rst), .QN(
        \cache[4][3][TAG][5] ) );
  DFFS_X1 \cache_reg[4][3][TAG][4]  ( .D(n253), .CK(net19313), .SN(rst), .QN(
        \cache[4][3][TAG][4] ) );
  DFFS_X1 \cache_reg[4][3][TAG][3]  ( .D(n254), .CK(net19313), .SN(rst), .QN(
        \cache[4][3][TAG][3] ) );
  DFFS_X1 \cache_reg[4][3][TAG][2]  ( .D(n255), .CK(net19313), .SN(rst), .QN(
        \cache[4][3][TAG][2] ) );
  DFFS_X1 \cache_reg[4][3][TAG][1]  ( .D(n256), .CK(net19313), .SN(rst), .QN(
        \cache[4][3][TAG][1] ) );
  DFFS_X1 \cache_reg[4][3][TAG][0]  ( .D(n257), .CK(net19313), .SN(rst), .QN(
        \cache[4][3][TAG][0] ) );
  DFFS_X1 \cache_reg[5][3][TAG][7]  ( .D(n250), .CK(net19373), .SN(rst), .QN(
        \cache[5][3][TAG][7] ) );
  DFFS_X1 \cache_reg[5][3][TAG][6]  ( .D(n251), .CK(net19373), .SN(rst), .QN(
        \cache[5][3][TAG][6] ) );
  DFFS_X1 \cache_reg[5][3][TAG][5]  ( .D(n252), .CK(net19373), .SN(rst), .QN(
        \cache[5][3][TAG][5] ) );
  DFFS_X1 \cache_reg[5][3][TAG][4]  ( .D(n253), .CK(net19373), .SN(rst), .QN(
        \cache[5][3][TAG][4] ) );
  DFFS_X1 \cache_reg[5][3][TAG][3]  ( .D(n254), .CK(net19373), .SN(rst), .QN(
        \cache[5][3][TAG][3] ) );
  DFFS_X1 \cache_reg[5][3][TAG][2]  ( .D(n255), .CK(net19373), .SN(rst), .QN(
        \cache[5][3][TAG][2] ) );
  DFFS_X1 \cache_reg[5][3][TAG][1]  ( .D(n256), .CK(net19373), .SN(rst), .QN(
        \cache[5][3][TAG][1] ) );
  DFFS_X1 \cache_reg[5][3][TAG][0]  ( .D(n257), .CK(net19373), .SN(rst), .QN(
        \cache[5][3][TAG][0] ) );
  DFFS_X1 \cache_reg[6][3][TAG][7]  ( .D(n250), .CK(net19433), .SN(rst), .QN(
        \cache[6][3][TAG][7] ) );
  DFFS_X1 \cache_reg[6][3][TAG][6]  ( .D(n251), .CK(net19433), .SN(rst), .QN(
        \cache[6][3][TAG][6] ) );
  DFFS_X1 \cache_reg[6][3][TAG][5]  ( .D(n252), .CK(net19433), .SN(rst), .QN(
        \cache[6][3][TAG][5] ) );
  DFFS_X1 \cache_reg[6][3][TAG][4]  ( .D(n253), .CK(net19433), .SN(rst), .QN(
        \cache[6][3][TAG][4] ) );
  DFFS_X1 \cache_reg[6][3][TAG][3]  ( .D(n254), .CK(net19433), .SN(rst), .QN(
        \cache[6][3][TAG][3] ) );
  DFFS_X1 \cache_reg[6][3][TAG][2]  ( .D(n255), .CK(net19433), .SN(rst), .QN(
        \cache[6][3][TAG][2] ) );
  DFFS_X1 \cache_reg[6][3][TAG][1]  ( .D(n256), .CK(net19433), .SN(rst), .QN(
        \cache[6][3][TAG][1] ) );
  DFFS_X1 \cache_reg[6][3][TAG][0]  ( .D(n257), .CK(net19433), .SN(rst), .QN(
        \cache[6][3][TAG][0] ) );
  DFFS_X1 \cache_reg[7][3][TAG][7]  ( .D(n250), .CK(net19493), .SN(rst), .QN(
        \cache[7][3][TAG][7] ) );
  DFFS_X1 \cache_reg[7][3][TAG][6]  ( .D(n251), .CK(net19493), .SN(rst), .QN(
        \cache[7][3][TAG][6] ) );
  DFFS_X1 \cache_reg[7][3][TAG][5]  ( .D(n252), .CK(net19493), .SN(rst), .QN(
        \cache[7][3][TAG][5] ) );
  DFFS_X1 \cache_reg[7][3][TAG][4]  ( .D(n253), .CK(net19493), .SN(rst), .QN(
        \cache[7][3][TAG][4] ) );
  DFFS_X1 \cache_reg[7][3][TAG][3]  ( .D(n254), .CK(net19493), .SN(rst), .QN(
        \cache[7][3][TAG][3] ) );
  DFFS_X1 \cache_reg[7][3][TAG][2]  ( .D(n255), .CK(net19493), .SN(rst), .QN(
        \cache[7][3][TAG][2] ) );
  DFFS_X1 \cache_reg[7][3][TAG][1]  ( .D(n256), .CK(net19493), .SN(rst), .QN(
        \cache[7][3][TAG][1] ) );
  DFFS_X1 \cache_reg[7][3][TAG][0]  ( .D(n257), .CK(net19493), .SN(rst), .QN(
        \cache[7][3][TAG][0] ) );
  DFFS_X1 \cache_reg[7][1][YOUTH][2]  ( .D(N2819), .CK(net19473), .SN(rst), 
        .Q(\cache[7][1][YOUTH][2] ) );
  DFFS_X1 \cache_reg[6][1][YOUTH][2]  ( .D(N2843), .CK(net19413), .SN(rst), 
        .Q(\cache[6][1][YOUTH][2] ) );
  DFFS_X1 \cache_reg[5][1][YOUTH][2]  ( .D(N2867), .CK(net19353), .SN(rst), 
        .Q(\cache[5][1][YOUTH][2] ) );
  DFFS_X1 \cache_reg[4][1][YOUTH][2]  ( .D(N2891), .CK(net19293), .SN(rst), 
        .Q(\cache[4][1][YOUTH][2] ) );
  DFFS_X1 \cache_reg[3][1][YOUTH][2]  ( .D(N2915), .CK(net19233), .SN(rst), 
        .Q(\cache[3][1][YOUTH][2] ) );
  DFFS_X1 \cache_reg[2][1][YOUTH][2]  ( .D(N2939), .CK(net19173), .SN(rst), 
        .Q(\cache[2][1][YOUTH][2] ) );
  DFFS_X1 \cache_reg[1][1][YOUTH][2]  ( .D(N2963), .CK(net19113), .SN(rst), 
        .Q(\cache[1][1][YOUTH][2] ) );
  DFFS_X1 \cache_reg[0][1][YOUTH][2]  ( .D(N2987), .CK(net19053), .SN(rst), 
        .Q(\cache[0][1][YOUTH][2] ) );
  DFFS_X1 \cache_reg[7][0][YOUTH][0]  ( .D(N2823), .CK(net19458), .SN(rst), 
        .Q(\cache[7][0][YOUTH][0] ) );
  DFFS_X1 \last_hit_index_reg[1]  ( .D(\hit_index[1] ), .CK(net19518), .SN(rst), .Q(\last_hit_index[1] ), .QN(n120) );
  DFFS_X1 \cache_reg[0][2][YOUTH][2]  ( .D(N2981), .CK(net19068), .SN(rst), 
        .Q(\cache[0][2][YOUTH][2] ) );
  DFFS_X1 \cache_reg[0][2][YOUTH][1]  ( .D(N2980), .CK(net19068), .SN(rst), 
        .Q(\cache[0][2][YOUTH][1] ) );
  DFFS_X1 \cache_reg[0][2][YOUTH][0]  ( .D(N2979), .CK(net19068), .SN(rst), 
        .Q(\cache[0][2][YOUTH][0] ) );
  DFFS_X1 \cache_reg[1][2][YOUTH][2]  ( .D(N2957), .CK(net19128), .SN(rst), 
        .Q(\cache[1][2][YOUTH][2] ) );
  DFFS_X1 \cache_reg[1][2][YOUTH][1]  ( .D(N2956), .CK(net19128), .SN(rst), 
        .Q(\cache[1][2][YOUTH][1] ) );
  DFFS_X1 \cache_reg[1][2][YOUTH][0]  ( .D(N2955), .CK(net19128), .SN(rst), 
        .Q(\cache[1][2][YOUTH][0] ) );
  DFFS_X1 \cache_reg[2][2][YOUTH][2]  ( .D(N2933), .CK(net19188), .SN(rst), 
        .Q(\cache[2][2][YOUTH][2] ) );
  DFFS_X1 \cache_reg[2][2][YOUTH][1]  ( .D(N2932), .CK(net19188), .SN(rst), 
        .Q(\cache[2][2][YOUTH][1] ) );
  DFFS_X1 \cache_reg[2][2][YOUTH][0]  ( .D(N2931), .CK(net19188), .SN(rst), 
        .Q(\cache[2][2][YOUTH][0] ) );
  DFFS_X1 \cache_reg[3][2][YOUTH][2]  ( .D(N2909), .CK(net19248), .SN(rst), 
        .Q(\cache[3][2][YOUTH][2] ) );
  DFFS_X1 \cache_reg[3][2][YOUTH][1]  ( .D(N2908), .CK(net19248), .SN(rst), 
        .Q(\cache[3][2][YOUTH][1] ) );
  DFFS_X1 \cache_reg[3][2][YOUTH][0]  ( .D(N2907), .CK(net19248), .SN(rst), 
        .Q(\cache[3][2][YOUTH][0] ) );
  DFFS_X1 \cache_reg[4][2][YOUTH][2]  ( .D(N2885), .CK(net19308), .SN(rst), 
        .Q(\cache[4][2][YOUTH][2] ) );
  DFFS_X1 \cache_reg[4][2][YOUTH][1]  ( .D(N2884), .CK(net19308), .SN(rst), 
        .Q(\cache[4][2][YOUTH][1] ) );
  DFFS_X1 \cache_reg[4][2][YOUTH][0]  ( .D(N2883), .CK(net19308), .SN(rst), 
        .Q(\cache[4][2][YOUTH][0] ) );
  DFFS_X1 \cache_reg[5][2][YOUTH][2]  ( .D(N2861), .CK(net19368), .SN(rst), 
        .Q(\cache[5][2][YOUTH][2] ) );
  DFFS_X1 \cache_reg[5][2][YOUTH][1]  ( .D(N2860), .CK(net19368), .SN(rst), 
        .Q(\cache[5][2][YOUTH][1] ) );
  DFFS_X1 \cache_reg[5][2][YOUTH][0]  ( .D(N2859), .CK(net19368), .SN(rst), 
        .Q(\cache[5][2][YOUTH][0] ) );
  DFFS_X1 \cache_reg[6][2][YOUTH][2]  ( .D(N2837), .CK(net19428), .SN(rst), 
        .Q(\cache[6][2][YOUTH][2] ) );
  DFFS_X1 \cache_reg[6][2][YOUTH][1]  ( .D(N2836), .CK(net19428), .SN(rst), 
        .Q(\cache[6][2][YOUTH][1] ) );
  DFFS_X1 \cache_reg[6][2][YOUTH][0]  ( .D(N2835), .CK(net19428), .SN(rst), 
        .Q(\cache[6][2][YOUTH][0] ) );
  DFFS_X1 \cache_reg[7][2][YOUTH][2]  ( .D(N2813), .CK(net19488), .SN(rst), 
        .Q(\cache[7][2][YOUTH][2] ) );
  DFFS_X1 \cache_reg[7][2][YOUTH][1]  ( .D(N2812), .CK(net19488), .SN(rst), 
        .Q(\cache[7][2][YOUTH][1] ) );
  DFFS_X1 \cache_reg[7][2][YOUTH][0]  ( .D(N2811), .CK(net19488), .SN(rst), 
        .Q(\cache[7][2][YOUTH][0] ) );
  DFFS_X1 \cache_reg[7][0][YOUTH][2]  ( .D(N2825), .CK(net19458), .SN(rst), 
        .Q(\cache[7][0][YOUTH][2] ) );
  DFFS_X1 \cache_reg[6][0][YOUTH][2]  ( .D(N2849), .CK(net19398), .SN(rst), 
        .Q(\cache[6][0][YOUTH][2] ) );
  DFFS_X1 \cache_reg[5][0][YOUTH][2]  ( .D(N2873), .CK(net19338), .SN(rst), 
        .Q(\cache[5][0][YOUTH][2] ) );
  DFFS_X1 \cache_reg[4][0][YOUTH][2]  ( .D(N2897), .CK(net19278), .SN(rst), 
        .Q(\cache[4][0][YOUTH][2] ) );
  DFFS_X1 \cache_reg[3][0][YOUTH][2]  ( .D(N2921), .CK(net19218), .SN(rst), 
        .Q(\cache[3][0][YOUTH][2] ) );
  DFFS_X1 \cache_reg[2][0][YOUTH][2]  ( .D(N2945), .CK(net19158), .SN(rst), 
        .Q(\cache[2][0][YOUTH][2] ) );
  DFFS_X1 \cache_reg[1][0][YOUTH][2]  ( .D(N2969), .CK(net19098), .SN(rst), 
        .Q(\cache[1][0][YOUTH][2] ) );
  DFFS_X1 \cache_reg[0][0][YOUTH][2]  ( .D(N2993), .CK(net19038), .SN(rst), 
        .Q(\cache[0][0][YOUTH][2] ) );
  DFFS_X1 \cache_reg[0][0][YOUTH][1]  ( .D(N2992), .CK(net19038), .SN(rst), 
        .Q(\cache[0][0][YOUTH][1] ) );
  DFFS_X1 \cache_reg[0][0][YOUTH][0]  ( .D(N2991), .CK(net19038), .SN(rst), 
        .Q(\cache[0][0][YOUTH][0] ) );
  DFFS_X1 \cache_reg[1][0][YOUTH][1]  ( .D(N2968), .CK(net19098), .SN(rst), 
        .Q(\cache[1][0][YOUTH][1] ) );
  DFFS_X1 \cache_reg[1][0][YOUTH][0]  ( .D(N2967), .CK(net19098), .SN(rst), 
        .Q(\cache[1][0][YOUTH][0] ) );
  DFFS_X1 \cache_reg[2][0][YOUTH][1]  ( .D(N2944), .CK(net19158), .SN(rst), 
        .Q(\cache[2][0][YOUTH][1] ) );
  DFFS_X1 \cache_reg[2][0][YOUTH][0]  ( .D(N2943), .CK(net19158), .SN(rst), 
        .Q(\cache[2][0][YOUTH][0] ) );
  DFFS_X1 \cache_reg[3][0][YOUTH][1]  ( .D(N2920), .CK(net19218), .SN(rst), 
        .Q(\cache[3][0][YOUTH][1] ) );
  DFFS_X1 \cache_reg[3][0][YOUTH][0]  ( .D(N2919), .CK(net19218), .SN(rst), 
        .Q(\cache[3][0][YOUTH][0] ) );
  DFFS_X1 \cache_reg[4][0][YOUTH][1]  ( .D(N2896), .CK(net19278), .SN(rst), 
        .Q(\cache[4][0][YOUTH][1] ) );
  DFFS_X1 \cache_reg[4][0][YOUTH][0]  ( .D(N2895), .CK(net19278), .SN(rst), 
        .Q(\cache[4][0][YOUTH][0] ) );
  DFFS_X1 \cache_reg[5][0][YOUTH][1]  ( .D(N2872), .CK(net19338), .SN(rst), 
        .Q(\cache[5][0][YOUTH][1] ) );
  DFFS_X1 \cache_reg[5][0][YOUTH][0]  ( .D(N2871), .CK(net19338), .SN(rst), 
        .Q(\cache[5][0][YOUTH][0] ) );
  DFFS_X1 \cache_reg[6][0][YOUTH][1]  ( .D(N2848), .CK(net19398), .SN(rst), 
        .Q(\cache[6][0][YOUTH][1] ) );
  DFFS_X1 \cache_reg[6][0][YOUTH][0]  ( .D(N2847), .CK(net19398), .SN(rst), 
        .Q(\cache[6][0][YOUTH][0] ) );
  DFFS_X1 \cache_reg[7][0][YOUTH][1]  ( .D(N2824), .CK(net19458), .SN(rst), 
        .Q(\cache[7][0][YOUTH][1] ) );
  DFFS_X1 \cache_reg[0][3][YOUTH][1]  ( .D(N2974), .CK(net19083), .SN(rst), 
        .Q(\cache[0][3][YOUTH][1] ) );
  DFFS_X1 \cache_reg[1][3][YOUTH][1]  ( .D(N2950), .CK(net19143), .SN(rst), 
        .Q(\cache[1][3][YOUTH][1] ) );
  DFFS_X1 \cache_reg[1][3][YOUTH][0]  ( .D(N2949), .CK(net19143), .SN(rst), 
        .Q(\cache[1][3][YOUTH][0] ) );
  DFFS_X1 \cache_reg[2][3][YOUTH][1]  ( .D(N2926), .CK(net19203), .SN(rst), 
        .Q(\cache[2][3][YOUTH][1] ) );
  DFFS_X1 \cache_reg[2][3][YOUTH][0]  ( .D(N2925), .CK(net19203), .SN(rst), 
        .Q(\cache[2][3][YOUTH][0] ) );
  DFFS_X1 \cache_reg[3][3][YOUTH][1]  ( .D(N2902), .CK(net19263), .SN(rst), 
        .Q(\cache[3][3][YOUTH][1] ) );
  DFFS_X1 \cache_reg[3][3][YOUTH][0]  ( .D(N2901), .CK(net19263), .SN(rst), 
        .Q(\cache[3][3][YOUTH][0] ) );
  DFFS_X1 \cache_reg[4][3][YOUTH][1]  ( .D(N2878), .CK(net19323), .SN(rst), 
        .Q(\cache[4][3][YOUTH][1] ) );
  DFFS_X1 \cache_reg[4][3][YOUTH][0]  ( .D(N2877), .CK(net19323), .SN(rst), 
        .Q(\cache[4][3][YOUTH][0] ) );
  DFFS_X1 \cache_reg[5][3][YOUTH][1]  ( .D(N2854), .CK(net19383), .SN(rst), 
        .Q(\cache[5][3][YOUTH][1] ) );
  DFFS_X1 \cache_reg[5][3][YOUTH][0]  ( .D(N2853), .CK(net19383), .SN(rst), 
        .Q(\cache[5][3][YOUTH][0] ) );
  DFFS_X1 \cache_reg[6][3][YOUTH][1]  ( .D(N2830), .CK(net19443), .SN(rst), 
        .Q(\cache[6][3][YOUTH][1] ) );
  DFFS_X1 \cache_reg[6][3][YOUTH][0]  ( .D(N2829), .CK(net19443), .SN(rst), 
        .Q(\cache[6][3][YOUTH][0] ) );
  DFFS_X1 \cache_reg[7][3][YOUTH][1]  ( .D(N2806), .CK(net19503), .SN(rst), 
        .Q(\cache[7][3][YOUTH][1] ) );
  DFFS_X1 \cache_reg[7][3][YOUTH][0]  ( .D(N2805), .CK(net19503), .SN(rst), 
        .Q(\cache[7][3][YOUTH][0] ) );
  DFFS_X1 \cache_reg[7][3][YOUTH][2]  ( .D(N2807), .CK(net19503), .SN(rst), 
        .Q(\cache[7][3][YOUTH][2] ) );
  DFFS_X1 \cache_reg[6][3][YOUTH][2]  ( .D(N2831), .CK(net19443), .SN(rst), 
        .Q(\cache[6][3][YOUTH][2] ) );
  DFFS_X1 \cache_reg[5][3][YOUTH][2]  ( .D(N2855), .CK(net19383), .SN(rst), 
        .Q(\cache[5][3][YOUTH][2] ) );
  DFFS_X1 \cache_reg[4][3][YOUTH][2]  ( .D(N2879), .CK(net19323), .SN(rst), 
        .Q(\cache[4][3][YOUTH][2] ) );
  DFFS_X1 \cache_reg[3][3][YOUTH][2]  ( .D(N2903), .CK(net19263), .SN(rst), 
        .Q(\cache[3][3][YOUTH][2] ) );
  DFFS_X1 \cache_reg[2][3][YOUTH][2]  ( .D(N2927), .CK(net19203), .SN(rst), 
        .Q(\cache[2][3][YOUTH][2] ) );
  DFFS_X1 \cache_reg[1][3][YOUTH][2]  ( .D(N2951), .CK(net19143), .SN(rst), 
        .Q(\cache[1][3][YOUTH][2] ) );
  DFFS_X1 \cache_reg[0][3][YOUTH][2]  ( .D(N2975), .CK(net19083), .SN(rst), 
        .Q(\cache[0][3][YOUTH][2] ) );
  DFFR_X1 \cache_reg[0][0][DATA][29]  ( .D(n300), .CK(net19033), .RN(rst), .Q(
        \cache[0][0][DATA][29] ) );
  DFFR_X1 \cache_reg[0][0][DATA][28]  ( .D(n298), .CK(net19033), .RN(rst), .Q(
        \cache[0][0][DATA][28] ) );
  DFFR_X1 \cache_reg[0][0][DATA][27]  ( .D(n296), .CK(net19033), .RN(rst), .Q(
        \cache[0][0][DATA][27] ) );
  DFFR_X1 \cache_reg[0][0][DATA][26]  ( .D(n294), .CK(net19033), .RN(rst), .Q(
        \cache[0][0][DATA][26] ) );
  DFFR_X1 \cache_reg[0][0][DATA][25]  ( .D(n292), .CK(net19033), .RN(rst), .Q(
        \cache[0][0][DATA][25] ) );
  DFFR_X1 \cache_reg[0][0][DATA][24]  ( .D(n290), .CK(net19033), .RN(rst), .Q(
        \cache[0][0][DATA][24] ) );
  DFFR_X1 \cache_reg[0][0][DATA][23]  ( .D(n288), .CK(net19033), .RN(rst), .Q(
        \cache[0][0][DATA][23] ) );
  DFFR_X1 \cache_reg[0][0][DATA][22]  ( .D(n286), .CK(net19033), .RN(rst), .Q(
        \cache[0][0][DATA][22] ) );
  DFFR_X1 \cache_reg[0][0][DATA][21]  ( .D(n44), .CK(net19033), .RN(rst), .Q(
        \cache[0][0][DATA][21] ) );
  DFFR_X1 \cache_reg[0][0][DATA][20]  ( .D(n42), .CK(net19033), .RN(rst), .Q(
        \cache[0][0][DATA][20] ) );
  DFFR_X1 \cache_reg[0][0][DATA][19]  ( .D(n48), .CK(net19033), .RN(rst), .Q(
        \cache[0][0][DATA][19] ) );
  DFFR_X1 \cache_reg[0][0][DATA][18]  ( .D(n46), .CK(net19033), .RN(rst), .Q(
        \cache[0][0][DATA][18] ) );
  DFFR_X1 \cache_reg[0][0][DATA][17]  ( .D(n47), .CK(net19033), .RN(rst), .Q(
        \cache[0][0][DATA][17] ) );
  DFFR_X1 \cache_reg[0][0][DATA][16]  ( .D(n279), .CK(net19033), .RN(rst), .Q(
        \cache[0][0][DATA][16] ) );
  DFFR_X1 \cache_reg[0][0][DATA][15]  ( .D(n45), .CK(net19033), .RN(rst), .Q(
        \cache[0][0][DATA][15] ) );
  DFFR_X1 \cache_reg[0][0][DATA][14]  ( .D(n35), .CK(net19033), .RN(rst), .Q(
        \cache[0][0][DATA][14] ) );
  DFFR_X1 \cache_reg[0][0][DATA][13]  ( .D(n52), .CK(net19033), .RN(rst), .Q(
        \cache[0][0][DATA][13] ) );
  DFFR_X1 \cache_reg[0][0][DATA][12]  ( .D(n50), .CK(net19033), .RN(rst), .Q(
        \cache[0][0][DATA][12] ) );
  DFFR_X1 \cache_reg[0][0][DATA][11]  ( .D(n51), .CK(net19033), .RN(rst), .Q(
        \cache[0][0][DATA][11] ) );
  DFFR_X1 \cache_reg[0][0][DATA][10]  ( .D(n49), .CK(net19033), .RN(rst), .Q(
        \cache[0][0][DATA][10] ) );
  DFFR_X1 \cache_reg[0][0][DATA][9]  ( .D(n43), .CK(net19033), .RN(rst), .Q(
        \cache[0][0][DATA][9] ) );
  DFFR_X1 \cache_reg[0][0][DATA][8]  ( .D(n270), .CK(net19033), .RN(rst), .Q(
        \cache[0][0][DATA][8] ) );
  DFFR_X1 \cache_reg[0][0][DATA][7]  ( .D(n204), .CK(net19033), .RN(rst), .Q(
        \cache[0][0][DATA][7] ) );
  DFFR_X1 \cache_reg[0][0][DATA][6]  ( .D(n222), .CK(net19033), .RN(rst), .Q(
        \cache[0][0][DATA][6] ) );
  DFFR_X1 \cache_reg[0][0][DATA][5]  ( .D(n266), .CK(net19033), .RN(rst), .Q(
        \cache[0][0][DATA][5] ) );
  DFFR_X1 \cache_reg[0][0][DATA][4]  ( .D(n264), .CK(net19033), .RN(rst), .Q(
        \cache[0][0][DATA][4] ) );
  DFFR_X1 \cache_reg[0][0][DATA][3]  ( .D(n262), .CK(net19033), .RN(rst), .Q(
        \cache[0][0][DATA][3] ) );
  DFFR_X1 \cache_reg[0][0][DATA][2]  ( .D(n260), .CK(net19033), .RN(rst), .Q(
        \cache[0][0][DATA][2] ) );
  DFFR_X1 \cache_reg[0][0][DATA][1]  ( .D(n216), .CK(net19033), .RN(rst), .Q(
        \cache[0][0][DATA][1] ) );
  DFFR_X1 \cache_reg[0][0][DATA][0]  ( .D(n212), .CK(net19033), .RN(rst), .Q(
        \cache[0][0][DATA][0] ) );
  DFFR_X1 \cache_reg[1][0][DATA][29]  ( .D(n300), .CK(net19093), .RN(rst), .Q(
        \cache[1][0][DATA][29] ) );
  DFFR_X1 \cache_reg[1][0][DATA][28]  ( .D(n298), .CK(net19093), .RN(rst), .Q(
        \cache[1][0][DATA][28] ) );
  DFFR_X1 \cache_reg[1][0][DATA][27]  ( .D(n296), .CK(net19093), .RN(rst), .Q(
        \cache[1][0][DATA][27] ) );
  DFFR_X1 \cache_reg[1][0][DATA][26]  ( .D(n294), .CK(net19093), .RN(rst), .Q(
        \cache[1][0][DATA][26] ) );
  DFFR_X1 \cache_reg[1][0][DATA][25]  ( .D(n292), .CK(net19093), .RN(rst), .Q(
        \cache[1][0][DATA][25] ) );
  DFFR_X1 \cache_reg[1][0][DATA][24]  ( .D(n290), .CK(net19093), .RN(rst), .Q(
        \cache[1][0][DATA][24] ) );
  DFFR_X1 \cache_reg[1][0][DATA][23]  ( .D(n288), .CK(net19093), .RN(rst), .Q(
        \cache[1][0][DATA][23] ) );
  DFFR_X1 \cache_reg[1][0][DATA][22]  ( .D(n286), .CK(net19093), .RN(rst), .Q(
        \cache[1][0][DATA][22] ) );
  DFFR_X1 \cache_reg[1][0][DATA][21]  ( .D(n44), .CK(net19093), .RN(rst), .Q(
        \cache[1][0][DATA][21] ) );
  DFFR_X1 \cache_reg[1][0][DATA][20]  ( .D(n42), .CK(net19093), .RN(rst), .Q(
        \cache[1][0][DATA][20] ) );
  DFFR_X1 \cache_reg[1][0][DATA][19]  ( .D(n48), .CK(net19093), .RN(rst), .Q(
        \cache[1][0][DATA][19] ) );
  DFFR_X1 \cache_reg[1][0][DATA][18]  ( .D(n46), .CK(net19093), .RN(rst), .Q(
        \cache[1][0][DATA][18] ) );
  DFFR_X1 \cache_reg[1][0][DATA][17]  ( .D(n47), .CK(net19093), .RN(rst), .Q(
        \cache[1][0][DATA][17] ) );
  DFFR_X1 \cache_reg[1][0][DATA][16]  ( .D(n279), .CK(net19093), .RN(rst), .Q(
        \cache[1][0][DATA][16] ) );
  DFFR_X1 \cache_reg[1][0][DATA][15]  ( .D(n45), .CK(net19093), .RN(rst), .Q(
        \cache[1][0][DATA][15] ) );
  DFFR_X1 \cache_reg[1][0][DATA][14]  ( .D(n35), .CK(net19093), .RN(rst), .Q(
        \cache[1][0][DATA][14] ) );
  DFFR_X1 \cache_reg[1][0][DATA][13]  ( .D(n52), .CK(net19093), .RN(rst), .Q(
        \cache[1][0][DATA][13] ) );
  DFFR_X1 \cache_reg[1][0][DATA][12]  ( .D(n50), .CK(net19093), .RN(rst), .Q(
        \cache[1][0][DATA][12] ) );
  DFFR_X1 \cache_reg[1][0][DATA][11]  ( .D(n51), .CK(net19093), .RN(rst), .Q(
        \cache[1][0][DATA][11] ) );
  DFFR_X1 \cache_reg[1][0][DATA][10]  ( .D(n49), .CK(net19093), .RN(rst), .Q(
        \cache[1][0][DATA][10] ) );
  DFFR_X1 \cache_reg[1][0][DATA][9]  ( .D(n43), .CK(net19093), .RN(rst), .Q(
        \cache[1][0][DATA][9] ) );
  DFFR_X1 \cache_reg[1][0][DATA][8]  ( .D(n270), .CK(net19093), .RN(rst), .Q(
        \cache[1][0][DATA][8] ) );
  DFFR_X1 \cache_reg[1][0][DATA][7]  ( .D(n204), .CK(net19093), .RN(rst), .Q(
        \cache[1][0][DATA][7] ) );
  DFFR_X1 \cache_reg[1][0][DATA][6]  ( .D(n222), .CK(net19093), .RN(rst), .Q(
        \cache[1][0][DATA][6] ) );
  DFFR_X1 \cache_reg[1][0][DATA][5]  ( .D(n266), .CK(net19093), .RN(rst), .Q(
        \cache[1][0][DATA][5] ) );
  DFFR_X1 \cache_reg[1][0][DATA][4]  ( .D(n264), .CK(net19093), .RN(rst), .Q(
        \cache[1][0][DATA][4] ) );
  DFFR_X1 \cache_reg[1][0][DATA][3]  ( .D(n262), .CK(net19093), .RN(rst), .Q(
        \cache[1][0][DATA][3] ) );
  DFFR_X1 \cache_reg[1][0][DATA][2]  ( .D(n260), .CK(net19093), .RN(rst), .Q(
        \cache[1][0][DATA][2] ) );
  DFFR_X1 \cache_reg[1][0][DATA][1]  ( .D(n216), .CK(net19093), .RN(rst), .Q(
        \cache[1][0][DATA][1] ) );
  DFFR_X1 \cache_reg[1][0][DATA][0]  ( .D(n212), .CK(net19093), .RN(rst), .Q(
        \cache[1][0][DATA][0] ) );
  DFFR_X1 \cache_reg[2][0][DATA][29]  ( .D(n300), .CK(net19153), .RN(rst), .Q(
        \cache[2][0][DATA][29] ) );
  DFFR_X1 \cache_reg[2][0][DATA][28]  ( .D(n298), .CK(net19153), .RN(rst), .Q(
        \cache[2][0][DATA][28] ) );
  DFFR_X1 \cache_reg[2][0][DATA][27]  ( .D(n296), .CK(net19153), .RN(rst), .Q(
        \cache[2][0][DATA][27] ) );
  DFFR_X1 \cache_reg[2][0][DATA][26]  ( .D(n294), .CK(net19153), .RN(rst), .Q(
        \cache[2][0][DATA][26] ) );
  DFFR_X1 \cache_reg[2][0][DATA][25]  ( .D(n292), .CK(net19153), .RN(rst), .Q(
        \cache[2][0][DATA][25] ) );
  DFFR_X1 \cache_reg[2][0][DATA][24]  ( .D(n290), .CK(net19153), .RN(rst), .Q(
        \cache[2][0][DATA][24] ) );
  DFFR_X1 \cache_reg[2][0][DATA][23]  ( .D(n288), .CK(net19153), .RN(rst), .Q(
        \cache[2][0][DATA][23] ) );
  DFFR_X1 \cache_reg[2][0][DATA][22]  ( .D(n286), .CK(net19153), .RN(rst), .Q(
        \cache[2][0][DATA][22] ) );
  DFFR_X1 \cache_reg[2][0][DATA][21]  ( .D(n44), .CK(net19153), .RN(rst), .Q(
        \cache[2][0][DATA][21] ) );
  DFFR_X1 \cache_reg[2][0][DATA][20]  ( .D(n42), .CK(net19153), .RN(rst), .Q(
        \cache[2][0][DATA][20] ) );
  DFFR_X1 \cache_reg[2][0][DATA][19]  ( .D(n48), .CK(net19153), .RN(rst), .Q(
        \cache[2][0][DATA][19] ) );
  DFFR_X1 \cache_reg[2][0][DATA][18]  ( .D(n46), .CK(net19153), .RN(rst), .Q(
        \cache[2][0][DATA][18] ) );
  DFFR_X1 \cache_reg[2][0][DATA][17]  ( .D(n47), .CK(net19153), .RN(rst), .Q(
        \cache[2][0][DATA][17] ) );
  DFFR_X1 \cache_reg[2][0][DATA][16]  ( .D(n279), .CK(net19153), .RN(rst), .Q(
        \cache[2][0][DATA][16] ) );
  DFFR_X1 \cache_reg[2][0][DATA][15]  ( .D(n45), .CK(net19153), .RN(rst), .Q(
        \cache[2][0][DATA][15] ) );
  DFFR_X1 \cache_reg[2][0][DATA][14]  ( .D(n35), .CK(net19153), .RN(rst), .Q(
        \cache[2][0][DATA][14] ) );
  DFFR_X1 \cache_reg[2][0][DATA][13]  ( .D(n52), .CK(net19153), .RN(rst), .Q(
        \cache[2][0][DATA][13] ) );
  DFFR_X1 \cache_reg[2][0][DATA][12]  ( .D(n50), .CK(net19153), .RN(rst), .Q(
        \cache[2][0][DATA][12] ) );
  DFFR_X1 \cache_reg[2][0][DATA][11]  ( .D(n51), .CK(net19153), .RN(rst), .Q(
        \cache[2][0][DATA][11] ) );
  DFFR_X1 \cache_reg[2][0][DATA][10]  ( .D(n49), .CK(net19153), .RN(rst), .Q(
        \cache[2][0][DATA][10] ) );
  DFFR_X1 \cache_reg[2][0][DATA][9]  ( .D(n43), .CK(net19153), .RN(rst), .Q(
        \cache[2][0][DATA][9] ) );
  DFFR_X1 \cache_reg[2][0][DATA][8]  ( .D(n270), .CK(net19153), .RN(rst), .Q(
        \cache[2][0][DATA][8] ) );
  DFFR_X1 \cache_reg[2][0][DATA][7]  ( .D(n204), .CK(net19153), .RN(rst), .Q(
        \cache[2][0][DATA][7] ) );
  DFFR_X1 \cache_reg[2][0][DATA][6]  ( .D(n222), .CK(net19153), .RN(rst), .Q(
        \cache[2][0][DATA][6] ) );
  DFFR_X1 \cache_reg[2][0][DATA][5]  ( .D(n266), .CK(net19153), .RN(rst), .Q(
        \cache[2][0][DATA][5] ) );
  DFFR_X1 \cache_reg[2][0][DATA][4]  ( .D(n264), .CK(net19153), .RN(rst), .Q(
        \cache[2][0][DATA][4] ) );
  DFFR_X1 \cache_reg[2][0][DATA][3]  ( .D(n262), .CK(net19153), .RN(rst), .Q(
        \cache[2][0][DATA][3] ) );
  DFFR_X1 \cache_reg[2][0][DATA][2]  ( .D(n260), .CK(net19153), .RN(rst), .Q(
        \cache[2][0][DATA][2] ) );
  DFFR_X1 \cache_reg[2][0][DATA][1]  ( .D(n216), .CK(net19153), .RN(rst), .Q(
        \cache[2][0][DATA][1] ) );
  DFFR_X1 \cache_reg[2][0][DATA][0]  ( .D(n212), .CK(net19153), .RN(rst), .Q(
        \cache[2][0][DATA][0] ) );
  DFFR_X1 \cache_reg[3][0][DATA][29]  ( .D(n300), .CK(net19213), .RN(rst), .Q(
        \cache[3][0][DATA][29] ) );
  DFFR_X1 \cache_reg[3][0][DATA][28]  ( .D(n298), .CK(net19213), .RN(rst), .Q(
        \cache[3][0][DATA][28] ) );
  DFFR_X1 \cache_reg[3][0][DATA][27]  ( .D(n296), .CK(net19213), .RN(rst), .Q(
        \cache[3][0][DATA][27] ) );
  DFFR_X1 \cache_reg[3][0][DATA][26]  ( .D(n294), .CK(net19213), .RN(rst), .Q(
        \cache[3][0][DATA][26] ) );
  DFFR_X1 \cache_reg[3][0][DATA][25]  ( .D(n292), .CK(net19213), .RN(rst), .Q(
        \cache[3][0][DATA][25] ) );
  DFFR_X1 \cache_reg[3][0][DATA][24]  ( .D(n290), .CK(net19213), .RN(rst), .Q(
        \cache[3][0][DATA][24] ) );
  DFFR_X1 \cache_reg[3][0][DATA][23]  ( .D(n288), .CK(net19213), .RN(rst), .Q(
        \cache[3][0][DATA][23] ) );
  DFFR_X1 \cache_reg[3][0][DATA][22]  ( .D(n286), .CK(net19213), .RN(rst), .Q(
        \cache[3][0][DATA][22] ) );
  DFFR_X1 \cache_reg[3][0][DATA][21]  ( .D(n44), .CK(net19213), .RN(rst), .Q(
        \cache[3][0][DATA][21] ) );
  DFFR_X1 \cache_reg[3][0][DATA][20]  ( .D(n42), .CK(net19213), .RN(rst), .Q(
        \cache[3][0][DATA][20] ) );
  DFFR_X1 \cache_reg[3][0][DATA][19]  ( .D(n48), .CK(net19213), .RN(rst), .Q(
        \cache[3][0][DATA][19] ) );
  DFFR_X1 \cache_reg[3][0][DATA][18]  ( .D(n46), .CK(net19213), .RN(rst), .Q(
        \cache[3][0][DATA][18] ) );
  DFFR_X1 \cache_reg[3][0][DATA][17]  ( .D(n47), .CK(net19213), .RN(rst), .Q(
        \cache[3][0][DATA][17] ) );
  DFFR_X1 \cache_reg[3][0][DATA][16]  ( .D(n279), .CK(net19213), .RN(rst), .Q(
        \cache[3][0][DATA][16] ) );
  DFFR_X1 \cache_reg[3][0][DATA][15]  ( .D(n45), .CK(net19213), .RN(rst), .Q(
        \cache[3][0][DATA][15] ) );
  DFFR_X1 \cache_reg[3][0][DATA][14]  ( .D(n35), .CK(net19213), .RN(rst), .Q(
        \cache[3][0][DATA][14] ) );
  DFFR_X1 \cache_reg[3][0][DATA][13]  ( .D(n52), .CK(net19213), .RN(rst), .Q(
        \cache[3][0][DATA][13] ) );
  DFFR_X1 \cache_reg[3][0][DATA][12]  ( .D(n50), .CK(net19213), .RN(rst), .Q(
        \cache[3][0][DATA][12] ) );
  DFFR_X1 \cache_reg[3][0][DATA][11]  ( .D(n51), .CK(net19213), .RN(rst), .Q(
        \cache[3][0][DATA][11] ) );
  DFFR_X1 \cache_reg[3][0][DATA][10]  ( .D(n49), .CK(net19213), .RN(rst), .Q(
        \cache[3][0][DATA][10] ) );
  DFFR_X1 \cache_reg[3][0][DATA][9]  ( .D(n43), .CK(net19213), .RN(rst), .Q(
        \cache[3][0][DATA][9] ) );
  DFFR_X1 \cache_reg[3][0][DATA][8]  ( .D(n270), .CK(net19213), .RN(rst), .Q(
        \cache[3][0][DATA][8] ) );
  DFFR_X1 \cache_reg[3][0][DATA][7]  ( .D(n204), .CK(net19213), .RN(rst), .Q(
        \cache[3][0][DATA][7] ) );
  DFFR_X1 \cache_reg[3][0][DATA][6]  ( .D(n222), .CK(net19213), .RN(rst), .Q(
        \cache[3][0][DATA][6] ) );
  DFFR_X1 \cache_reg[3][0][DATA][5]  ( .D(n266), .CK(net19213), .RN(rst), .Q(
        \cache[3][0][DATA][5] ) );
  DFFR_X1 \cache_reg[3][0][DATA][4]  ( .D(n264), .CK(net19213), .RN(rst), .Q(
        \cache[3][0][DATA][4] ) );
  DFFR_X1 \cache_reg[3][0][DATA][3]  ( .D(n262), .CK(net19213), .RN(rst), .Q(
        \cache[3][0][DATA][3] ) );
  DFFR_X1 \cache_reg[3][0][DATA][2]  ( .D(n260), .CK(net19213), .RN(rst), .Q(
        \cache[3][0][DATA][2] ) );
  DFFR_X1 \cache_reg[3][0][DATA][1]  ( .D(n216), .CK(net19213), .RN(rst), .Q(
        \cache[3][0][DATA][1] ) );
  DFFR_X1 \cache_reg[3][0][DATA][0]  ( .D(n212), .CK(net19213), .RN(rst), .Q(
        \cache[3][0][DATA][0] ) );
  DFFR_X1 \cache_reg[4][0][DATA][29]  ( .D(n300), .CK(net19273), .RN(rst), .Q(
        \cache[4][0][DATA][29] ) );
  DFFR_X1 \cache_reg[4][0][DATA][28]  ( .D(n298), .CK(net19273), .RN(rst), .Q(
        \cache[4][0][DATA][28] ) );
  DFFR_X1 \cache_reg[4][0][DATA][27]  ( .D(n296), .CK(net19273), .RN(rst), .Q(
        \cache[4][0][DATA][27] ) );
  DFFR_X1 \cache_reg[4][0][DATA][26]  ( .D(n294), .CK(net19273), .RN(rst), .Q(
        \cache[4][0][DATA][26] ) );
  DFFR_X1 \cache_reg[4][0][DATA][25]  ( .D(n292), .CK(net19273), .RN(rst), .Q(
        \cache[4][0][DATA][25] ) );
  DFFR_X1 \cache_reg[4][0][DATA][24]  ( .D(n290), .CK(net19273), .RN(rst), .Q(
        \cache[4][0][DATA][24] ) );
  DFFR_X1 \cache_reg[4][0][DATA][23]  ( .D(n288), .CK(net19273), .RN(rst), .Q(
        \cache[4][0][DATA][23] ) );
  DFFR_X1 \cache_reg[4][0][DATA][22]  ( .D(n286), .CK(net19273), .RN(rst), .Q(
        \cache[4][0][DATA][22] ) );
  DFFR_X1 \cache_reg[4][0][DATA][21]  ( .D(n44), .CK(net19273), .RN(rst), .Q(
        \cache[4][0][DATA][21] ) );
  DFFR_X1 \cache_reg[4][0][DATA][20]  ( .D(n42), .CK(net19273), .RN(rst), .Q(
        \cache[4][0][DATA][20] ) );
  DFFR_X1 \cache_reg[4][0][DATA][19]  ( .D(n48), .CK(net19273), .RN(rst), .Q(
        \cache[4][0][DATA][19] ) );
  DFFR_X1 \cache_reg[4][0][DATA][18]  ( .D(n46), .CK(net19273), .RN(rst), .Q(
        \cache[4][0][DATA][18] ) );
  DFFR_X1 \cache_reg[4][0][DATA][17]  ( .D(n47), .CK(net19273), .RN(rst), .Q(
        \cache[4][0][DATA][17] ) );
  DFFR_X1 \cache_reg[4][0][DATA][16]  ( .D(n279), .CK(net19273), .RN(rst), .Q(
        \cache[4][0][DATA][16] ) );
  DFFR_X1 \cache_reg[4][0][DATA][15]  ( .D(n45), .CK(net19273), .RN(rst), .Q(
        \cache[4][0][DATA][15] ) );
  DFFR_X1 \cache_reg[4][0][DATA][14]  ( .D(n35), .CK(net19273), .RN(rst), .Q(
        \cache[4][0][DATA][14] ) );
  DFFR_X1 \cache_reg[4][0][DATA][13]  ( .D(n52), .CK(net19273), .RN(rst), .Q(
        \cache[4][0][DATA][13] ) );
  DFFR_X1 \cache_reg[4][0][DATA][12]  ( .D(n50), .CK(net19273), .RN(rst), .Q(
        \cache[4][0][DATA][12] ) );
  DFFR_X1 \cache_reg[4][0][DATA][11]  ( .D(n51), .CK(net19273), .RN(rst), .Q(
        \cache[4][0][DATA][11] ) );
  DFFR_X1 \cache_reg[4][0][DATA][10]  ( .D(n49), .CK(net19273), .RN(rst), .Q(
        \cache[4][0][DATA][10] ) );
  DFFR_X1 \cache_reg[4][0][DATA][9]  ( .D(n43), .CK(net19273), .RN(rst), .Q(
        \cache[4][0][DATA][9] ) );
  DFFR_X1 \cache_reg[4][0][DATA][8]  ( .D(n270), .CK(net19273), .RN(rst), .Q(
        \cache[4][0][DATA][8] ) );
  DFFR_X1 \cache_reg[4][0][DATA][7]  ( .D(n204), .CK(net19273), .RN(rst), .Q(
        \cache[4][0][DATA][7] ) );
  DFFR_X1 \cache_reg[4][0][DATA][6]  ( .D(n222), .CK(net19273), .RN(rst), .Q(
        \cache[4][0][DATA][6] ) );
  DFFR_X1 \cache_reg[4][0][DATA][5]  ( .D(n266), .CK(net19273), .RN(rst), .Q(
        \cache[4][0][DATA][5] ) );
  DFFR_X1 \cache_reg[4][0][DATA][4]  ( .D(n264), .CK(net19273), .RN(rst), .Q(
        \cache[4][0][DATA][4] ) );
  DFFR_X1 \cache_reg[4][0][DATA][3]  ( .D(n262), .CK(net19273), .RN(rst), .Q(
        \cache[4][0][DATA][3] ) );
  DFFR_X1 \cache_reg[4][0][DATA][2]  ( .D(n260), .CK(net19273), .RN(rst), .Q(
        \cache[4][0][DATA][2] ) );
  DFFR_X1 \cache_reg[4][0][DATA][1]  ( .D(n216), .CK(net19273), .RN(rst), .Q(
        \cache[4][0][DATA][1] ) );
  DFFR_X1 \cache_reg[4][0][DATA][0]  ( .D(n212), .CK(net19273), .RN(rst), .Q(
        \cache[4][0][DATA][0] ) );
  DFFR_X1 \cache_reg[5][0][DATA][29]  ( .D(n300), .CK(net19333), .RN(rst), .Q(
        \cache[5][0][DATA][29] ) );
  DFFR_X1 \cache_reg[5][0][DATA][28]  ( .D(n298), .CK(net19333), .RN(rst), .Q(
        \cache[5][0][DATA][28] ) );
  DFFR_X1 \cache_reg[5][0][DATA][27]  ( .D(n296), .CK(net19333), .RN(rst), .Q(
        \cache[5][0][DATA][27] ) );
  DFFR_X1 \cache_reg[5][0][DATA][26]  ( .D(n294), .CK(net19333), .RN(rst), .Q(
        \cache[5][0][DATA][26] ) );
  DFFR_X1 \cache_reg[5][0][DATA][25]  ( .D(n292), .CK(net19333), .RN(rst), .Q(
        \cache[5][0][DATA][25] ) );
  DFFR_X1 \cache_reg[5][0][DATA][24]  ( .D(n290), .CK(net19333), .RN(rst), .Q(
        \cache[5][0][DATA][24] ) );
  DFFR_X1 \cache_reg[5][0][DATA][23]  ( .D(n288), .CK(net19333), .RN(rst), .Q(
        \cache[5][0][DATA][23] ) );
  DFFR_X1 \cache_reg[5][0][DATA][22]  ( .D(n286), .CK(net19333), .RN(rst), .Q(
        \cache[5][0][DATA][22] ) );
  DFFR_X1 \cache_reg[5][0][DATA][21]  ( .D(n44), .CK(net19333), .RN(rst), .Q(
        \cache[5][0][DATA][21] ) );
  DFFR_X1 \cache_reg[5][0][DATA][20]  ( .D(n42), .CK(net19333), .RN(rst), .Q(
        \cache[5][0][DATA][20] ) );
  DFFR_X1 \cache_reg[5][0][DATA][19]  ( .D(n48), .CK(net19333), .RN(rst), .Q(
        \cache[5][0][DATA][19] ) );
  DFFR_X1 \cache_reg[5][0][DATA][18]  ( .D(n46), .CK(net19333), .RN(rst), .Q(
        \cache[5][0][DATA][18] ) );
  DFFR_X1 \cache_reg[5][0][DATA][17]  ( .D(n47), .CK(net19333), .RN(rst), .Q(
        \cache[5][0][DATA][17] ) );
  DFFR_X1 \cache_reg[5][0][DATA][16]  ( .D(n279), .CK(net19333), .RN(rst), .Q(
        \cache[5][0][DATA][16] ) );
  DFFR_X1 \cache_reg[5][0][DATA][15]  ( .D(n45), .CK(net19333), .RN(rst), .Q(
        \cache[5][0][DATA][15] ) );
  DFFR_X1 \cache_reg[5][0][DATA][14]  ( .D(n35), .CK(net19333), .RN(rst), .Q(
        \cache[5][0][DATA][14] ) );
  DFFR_X1 \cache_reg[5][0][DATA][13]  ( .D(n52), .CK(net19333), .RN(rst), .Q(
        \cache[5][0][DATA][13] ) );
  DFFR_X1 \cache_reg[5][0][DATA][12]  ( .D(n50), .CK(net19333), .RN(rst), .Q(
        \cache[5][0][DATA][12] ) );
  DFFR_X1 \cache_reg[5][0][DATA][11]  ( .D(n51), .CK(net19333), .RN(rst), .Q(
        \cache[5][0][DATA][11] ) );
  DFFR_X1 \cache_reg[5][0][DATA][10]  ( .D(n49), .CK(net19333), .RN(rst), .Q(
        \cache[5][0][DATA][10] ) );
  DFFR_X1 \cache_reg[5][0][DATA][9]  ( .D(n43), .CK(net19333), .RN(rst), .Q(
        \cache[5][0][DATA][9] ) );
  DFFR_X1 \cache_reg[5][0][DATA][8]  ( .D(n270), .CK(net19333), .RN(rst), .Q(
        \cache[5][0][DATA][8] ) );
  DFFR_X1 \cache_reg[5][0][DATA][7]  ( .D(n204), .CK(net19333), .RN(rst), .Q(
        \cache[5][0][DATA][7] ) );
  DFFR_X1 \cache_reg[5][0][DATA][6]  ( .D(n222), .CK(net19333), .RN(rst), .Q(
        \cache[5][0][DATA][6] ) );
  DFFR_X1 \cache_reg[5][0][DATA][5]  ( .D(n266), .CK(net19333), .RN(rst), .Q(
        \cache[5][0][DATA][5] ) );
  DFFR_X1 \cache_reg[5][0][DATA][4]  ( .D(n264), .CK(net19333), .RN(rst), .Q(
        \cache[5][0][DATA][4] ) );
  DFFR_X1 \cache_reg[5][0][DATA][3]  ( .D(n262), .CK(net19333), .RN(rst), .Q(
        \cache[5][0][DATA][3] ) );
  DFFR_X1 \cache_reg[5][0][DATA][2]  ( .D(n260), .CK(net19333), .RN(rst), .Q(
        \cache[5][0][DATA][2] ) );
  DFFR_X1 \cache_reg[5][0][DATA][1]  ( .D(n216), .CK(net19333), .RN(rst), .Q(
        \cache[5][0][DATA][1] ) );
  DFFR_X1 \cache_reg[5][0][DATA][0]  ( .D(n212), .CK(net19333), .RN(rst), .Q(
        \cache[5][0][DATA][0] ) );
  DFFR_X1 \cache_reg[6][0][DATA][29]  ( .D(n300), .CK(net19393), .RN(rst), .Q(
        \cache[6][0][DATA][29] ) );
  DFFR_X1 \cache_reg[6][0][DATA][28]  ( .D(n298), .CK(net19393), .RN(rst), .Q(
        \cache[6][0][DATA][28] ) );
  DFFR_X1 \cache_reg[6][0][DATA][27]  ( .D(n296), .CK(net19393), .RN(rst), .Q(
        \cache[6][0][DATA][27] ) );
  DFFR_X1 \cache_reg[6][0][DATA][26]  ( .D(n294), .CK(net19393), .RN(rst), .Q(
        \cache[6][0][DATA][26] ) );
  DFFR_X1 \cache_reg[6][0][DATA][25]  ( .D(n292), .CK(net19393), .RN(rst), .Q(
        \cache[6][0][DATA][25] ) );
  DFFR_X1 \cache_reg[6][0][DATA][24]  ( .D(n290), .CK(net19393), .RN(rst), .Q(
        \cache[6][0][DATA][24] ) );
  DFFR_X1 \cache_reg[6][0][DATA][23]  ( .D(n288), .CK(net19393), .RN(rst), .Q(
        \cache[6][0][DATA][23] ) );
  DFFR_X1 \cache_reg[6][0][DATA][22]  ( .D(n286), .CK(net19393), .RN(rst), .Q(
        \cache[6][0][DATA][22] ) );
  DFFR_X1 \cache_reg[6][0][DATA][21]  ( .D(n44), .CK(net19393), .RN(rst), .Q(
        \cache[6][0][DATA][21] ) );
  DFFR_X1 \cache_reg[6][0][DATA][20]  ( .D(n42), .CK(net19393), .RN(rst), .Q(
        \cache[6][0][DATA][20] ) );
  DFFR_X1 \cache_reg[6][0][DATA][19]  ( .D(n48), .CK(net19393), .RN(rst), .Q(
        \cache[6][0][DATA][19] ) );
  DFFR_X1 \cache_reg[6][0][DATA][18]  ( .D(n46), .CK(net19393), .RN(rst), .Q(
        \cache[6][0][DATA][18] ) );
  DFFR_X1 \cache_reg[6][0][DATA][17]  ( .D(n47), .CK(net19393), .RN(rst), .Q(
        \cache[6][0][DATA][17] ) );
  DFFR_X1 \cache_reg[6][0][DATA][16]  ( .D(n279), .CK(net19393), .RN(rst), .Q(
        \cache[6][0][DATA][16] ) );
  DFFR_X1 \cache_reg[6][0][DATA][15]  ( .D(n45), .CK(net19393), .RN(rst), .Q(
        \cache[6][0][DATA][15] ) );
  DFFR_X1 \cache_reg[6][0][DATA][14]  ( .D(n35), .CK(net19393), .RN(rst), .Q(
        \cache[6][0][DATA][14] ) );
  DFFR_X1 \cache_reg[6][0][DATA][13]  ( .D(n52), .CK(net19393), .RN(rst), .Q(
        \cache[6][0][DATA][13] ) );
  DFFR_X1 \cache_reg[6][0][DATA][12]  ( .D(n50), .CK(net19393), .RN(rst), .Q(
        \cache[6][0][DATA][12] ) );
  DFFR_X1 \cache_reg[6][0][DATA][11]  ( .D(n51), .CK(net19393), .RN(rst), .Q(
        \cache[6][0][DATA][11] ) );
  DFFR_X1 \cache_reg[6][0][DATA][10]  ( .D(n49), .CK(net19393), .RN(rst), .Q(
        \cache[6][0][DATA][10] ) );
  DFFR_X1 \cache_reg[6][0][DATA][9]  ( .D(n43), .CK(net19393), .RN(rst), .Q(
        \cache[6][0][DATA][9] ) );
  DFFR_X1 \cache_reg[6][0][DATA][8]  ( .D(n270), .CK(net19393), .RN(rst), .Q(
        \cache[6][0][DATA][8] ) );
  DFFR_X1 \cache_reg[6][0][DATA][7]  ( .D(n204), .CK(net19393), .RN(rst), .Q(
        \cache[6][0][DATA][7] ) );
  DFFR_X1 \cache_reg[6][0][DATA][6]  ( .D(n222), .CK(net19393), .RN(rst), .Q(
        \cache[6][0][DATA][6] ) );
  DFFR_X1 \cache_reg[6][0][DATA][5]  ( .D(n266), .CK(net19393), .RN(rst), .Q(
        \cache[6][0][DATA][5] ) );
  DFFR_X1 \cache_reg[6][0][DATA][4]  ( .D(n264), .CK(net19393), .RN(rst), .Q(
        \cache[6][0][DATA][4] ) );
  DFFR_X1 \cache_reg[6][0][DATA][3]  ( .D(n262), .CK(net19393), .RN(rst), .Q(
        \cache[6][0][DATA][3] ) );
  DFFR_X1 \cache_reg[6][0][DATA][2]  ( .D(n260), .CK(net19393), .RN(rst), .Q(
        \cache[6][0][DATA][2] ) );
  DFFR_X1 \cache_reg[6][0][DATA][1]  ( .D(n216), .CK(net19393), .RN(rst), .Q(
        \cache[6][0][DATA][1] ) );
  DFFR_X1 \cache_reg[6][0][DATA][0]  ( .D(n212), .CK(net19393), .RN(rst), .Q(
        \cache[6][0][DATA][0] ) );
  DFFR_X1 \cache_reg[7][0][DATA][29]  ( .D(n300), .CK(net19453), .RN(rst), .Q(
        \cache[7][0][DATA][29] ) );
  DFFR_X1 \cache_reg[7][0][DATA][28]  ( .D(n298), .CK(net19453), .RN(rst), .Q(
        \cache[7][0][DATA][28] ) );
  DFFR_X1 \cache_reg[7][0][DATA][27]  ( .D(n296), .CK(net19453), .RN(rst), .Q(
        \cache[7][0][DATA][27] ) );
  DFFR_X1 \cache_reg[7][0][DATA][26]  ( .D(n294), .CK(net19453), .RN(rst), .Q(
        \cache[7][0][DATA][26] ) );
  DFFR_X1 \cache_reg[7][0][DATA][25]  ( .D(n292), .CK(net19453), .RN(rst), .Q(
        \cache[7][0][DATA][25] ) );
  DFFR_X1 \cache_reg[7][0][DATA][24]  ( .D(n290), .CK(net19453), .RN(rst), .Q(
        \cache[7][0][DATA][24] ) );
  DFFR_X1 \cache_reg[7][0][DATA][23]  ( .D(n288), .CK(net19453), .RN(rst), .Q(
        \cache[7][0][DATA][23] ) );
  DFFR_X1 \cache_reg[7][0][DATA][22]  ( .D(n286), .CK(net19453), .RN(rst), .Q(
        \cache[7][0][DATA][22] ) );
  DFFR_X1 \cache_reg[7][0][DATA][21]  ( .D(n44), .CK(net19453), .RN(rst), .Q(
        \cache[7][0][DATA][21] ) );
  DFFR_X1 \cache_reg[7][0][DATA][20]  ( .D(n42), .CK(net19453), .RN(rst), .Q(
        \cache[7][0][DATA][20] ) );
  DFFR_X1 \cache_reg[7][0][DATA][19]  ( .D(n48), .CK(net19453), .RN(rst), .Q(
        \cache[7][0][DATA][19] ) );
  DFFR_X1 \cache_reg[7][0][DATA][18]  ( .D(n46), .CK(net19453), .RN(rst), .Q(
        \cache[7][0][DATA][18] ) );
  DFFR_X1 \cache_reg[7][0][DATA][17]  ( .D(n47), .CK(net19453), .RN(rst), .Q(
        \cache[7][0][DATA][17] ) );
  DFFR_X1 \cache_reg[7][0][DATA][16]  ( .D(n279), .CK(net19453), .RN(rst), .Q(
        \cache[7][0][DATA][16] ) );
  DFFR_X1 \cache_reg[7][0][DATA][15]  ( .D(n45), .CK(net19453), .RN(rst), .Q(
        \cache[7][0][DATA][15] ) );
  DFFR_X1 \cache_reg[7][0][DATA][14]  ( .D(n35), .CK(net19453), .RN(rst), .Q(
        \cache[7][0][DATA][14] ) );
  DFFR_X1 \cache_reg[7][0][DATA][13]  ( .D(n52), .CK(net19453), .RN(rst), .Q(
        \cache[7][0][DATA][13] ) );
  DFFR_X1 \cache_reg[7][0][DATA][12]  ( .D(n50), .CK(net19453), .RN(rst), .Q(
        \cache[7][0][DATA][12] ) );
  DFFR_X1 \cache_reg[7][0][DATA][11]  ( .D(n51), .CK(net19453), .RN(rst), .Q(
        \cache[7][0][DATA][11] ) );
  DFFR_X1 \cache_reg[7][0][DATA][10]  ( .D(n49), .CK(net19453), .RN(rst), .Q(
        \cache[7][0][DATA][10] ) );
  DFFR_X1 \cache_reg[7][0][DATA][9]  ( .D(n43), .CK(net19453), .RN(rst), .Q(
        \cache[7][0][DATA][9] ) );
  DFFR_X1 \cache_reg[7][0][DATA][8]  ( .D(n270), .CK(net19453), .RN(rst), .Q(
        \cache[7][0][DATA][8] ) );
  DFFR_X1 \cache_reg[7][0][DATA][7]  ( .D(n204), .CK(net19453), .RN(rst), .Q(
        \cache[7][0][DATA][7] ) );
  DFFR_X1 \cache_reg[7][0][DATA][6]  ( .D(n222), .CK(net19453), .RN(rst), .Q(
        \cache[7][0][DATA][6] ) );
  DFFR_X1 \cache_reg[7][0][DATA][5]  ( .D(n266), .CK(net19453), .RN(rst), .Q(
        \cache[7][0][DATA][5] ) );
  DFFR_X1 \cache_reg[7][0][DATA][4]  ( .D(n264), .CK(net19453), .RN(rst), .Q(
        \cache[7][0][DATA][4] ) );
  DFFR_X1 \cache_reg[7][0][DATA][3]  ( .D(n262), .CK(net19453), .RN(rst), .Q(
        \cache[7][0][DATA][3] ) );
  DFFR_X1 \cache_reg[7][0][DATA][2]  ( .D(n260), .CK(net19453), .RN(rst), .Q(
        \cache[7][0][DATA][2] ) );
  DFFR_X1 \cache_reg[7][0][DATA][1]  ( .D(n216), .CK(net19453), .RN(rst), .Q(
        \cache[7][0][DATA][1] ) );
  DFFR_X1 \cache_reg[7][0][DATA][0]  ( .D(n212), .CK(net19453), .RN(rst), .Q(
        \cache[7][0][DATA][0] ) );
  DFFR_X1 \cache_reg[0][1][DATA][29]  ( .D(n300), .CK(net19048), .RN(rst), .Q(
        \cache[0][1][DATA][29] ) );
  DFFR_X1 \cache_reg[0][1][DATA][28]  ( .D(n298), .CK(net19048), .RN(rst), .Q(
        \cache[0][1][DATA][28] ) );
  DFFR_X1 \cache_reg[0][1][DATA][27]  ( .D(n296), .CK(net19048), .RN(rst), .Q(
        \cache[0][1][DATA][27] ) );
  DFFR_X1 \cache_reg[0][1][DATA][26]  ( .D(n294), .CK(net19048), .RN(rst), .Q(
        \cache[0][1][DATA][26] ) );
  DFFR_X1 \cache_reg[0][1][DATA][25]  ( .D(n292), .CK(net19048), .RN(rst), .Q(
        \cache[0][1][DATA][25] ) );
  DFFR_X1 \cache_reg[0][1][DATA][24]  ( .D(n290), .CK(net19048), .RN(rst), .Q(
        \cache[0][1][DATA][24] ) );
  DFFR_X1 \cache_reg[0][1][DATA][23]  ( .D(n288), .CK(net19048), .RN(rst), .Q(
        \cache[0][1][DATA][23] ) );
  DFFR_X1 \cache_reg[0][1][DATA][22]  ( .D(n286), .CK(net19048), .RN(rst), .Q(
        \cache[0][1][DATA][22] ) );
  DFFR_X1 \cache_reg[0][1][DATA][21]  ( .D(n44), .CK(net19048), .RN(rst), .Q(
        \cache[0][1][DATA][21] ) );
  DFFR_X1 \cache_reg[0][1][DATA][20]  ( .D(n42), .CK(net19048), .RN(rst), .Q(
        \cache[0][1][DATA][20] ) );
  DFFR_X1 \cache_reg[0][1][DATA][19]  ( .D(n48), .CK(net19048), .RN(rst), .Q(
        \cache[0][1][DATA][19] ) );
  DFFR_X1 \cache_reg[0][1][DATA][18]  ( .D(n46), .CK(net19048), .RN(rst), .Q(
        \cache[0][1][DATA][18] ) );
  DFFR_X1 \cache_reg[0][1][DATA][17]  ( .D(n47), .CK(net19048), .RN(rst), .Q(
        \cache[0][1][DATA][17] ) );
  DFFR_X1 \cache_reg[0][1][DATA][16]  ( .D(n279), .CK(net19048), .RN(rst), .Q(
        \cache[0][1][DATA][16] ) );
  DFFR_X1 \cache_reg[0][1][DATA][15]  ( .D(n45), .CK(net19048), .RN(rst), .Q(
        \cache[0][1][DATA][15] ) );
  DFFR_X1 \cache_reg[0][1][DATA][14]  ( .D(n35), .CK(net19048), .RN(rst), .Q(
        \cache[0][1][DATA][14] ) );
  DFFR_X1 \cache_reg[0][1][DATA][13]  ( .D(n52), .CK(net19048), .RN(rst), .Q(
        \cache[0][1][DATA][13] ) );
  DFFR_X1 \cache_reg[0][1][DATA][12]  ( .D(n50), .CK(net19048), .RN(rst), .Q(
        \cache[0][1][DATA][12] ) );
  DFFR_X1 \cache_reg[0][1][DATA][11]  ( .D(n51), .CK(net19048), .RN(rst), .Q(
        \cache[0][1][DATA][11] ) );
  DFFR_X1 \cache_reg[0][1][DATA][10]  ( .D(n49), .CK(net19048), .RN(rst), .Q(
        \cache[0][1][DATA][10] ) );
  DFFR_X1 \cache_reg[0][1][DATA][9]  ( .D(n43), .CK(net19048), .RN(rst), .Q(
        \cache[0][1][DATA][9] ) );
  DFFR_X1 \cache_reg[0][1][DATA][8]  ( .D(n270), .CK(net19048), .RN(rst), .Q(
        \cache[0][1][DATA][8] ) );
  DFFR_X1 \cache_reg[0][1][DATA][7]  ( .D(n204), .CK(net19048), .RN(rst), .Q(
        \cache[0][1][DATA][7] ) );
  DFFR_X1 \cache_reg[0][1][DATA][6]  ( .D(n222), .CK(net19048), .RN(rst), .Q(
        \cache[0][1][DATA][6] ) );
  DFFR_X1 \cache_reg[0][1][DATA][5]  ( .D(n266), .CK(net19048), .RN(rst), .Q(
        \cache[0][1][DATA][5] ) );
  DFFR_X1 \cache_reg[0][1][DATA][4]  ( .D(n264), .CK(net19048), .RN(rst), .Q(
        \cache[0][1][DATA][4] ) );
  DFFR_X1 \cache_reg[0][1][DATA][3]  ( .D(n262), .CK(net19048), .RN(rst), .Q(
        \cache[0][1][DATA][3] ) );
  DFFR_X1 \cache_reg[0][1][DATA][2]  ( .D(n260), .CK(net19048), .RN(rst), .Q(
        \cache[0][1][DATA][2] ) );
  DFFR_X1 \cache_reg[0][1][DATA][1]  ( .D(n216), .CK(net19048), .RN(rst), .Q(
        \cache[0][1][DATA][1] ) );
  DFFR_X1 \cache_reg[0][1][DATA][0]  ( .D(n212), .CK(net19048), .RN(rst), .Q(
        \cache[0][1][DATA][0] ) );
  DFFR_X1 \cache_reg[1][1][DATA][29]  ( .D(n300), .CK(net19108), .RN(rst), .Q(
        \cache[1][1][DATA][29] ) );
  DFFR_X1 \cache_reg[1][1][DATA][28]  ( .D(n298), .CK(net19108), .RN(rst), .Q(
        \cache[1][1][DATA][28] ) );
  DFFR_X1 \cache_reg[1][1][DATA][27]  ( .D(n296), .CK(net19108), .RN(rst), .Q(
        \cache[1][1][DATA][27] ) );
  DFFR_X1 \cache_reg[1][1][DATA][26]  ( .D(n294), .CK(net19108), .RN(rst), .Q(
        \cache[1][1][DATA][26] ) );
  DFFR_X1 \cache_reg[1][1][DATA][25]  ( .D(n292), .CK(net19108), .RN(rst), .Q(
        \cache[1][1][DATA][25] ) );
  DFFR_X1 \cache_reg[1][1][DATA][24]  ( .D(n290), .CK(net19108), .RN(rst), .Q(
        \cache[1][1][DATA][24] ) );
  DFFR_X1 \cache_reg[1][1][DATA][23]  ( .D(n288), .CK(net19108), .RN(rst), .Q(
        \cache[1][1][DATA][23] ) );
  DFFR_X1 \cache_reg[1][1][DATA][22]  ( .D(n286), .CK(net19108), .RN(rst), .Q(
        \cache[1][1][DATA][22] ) );
  DFFR_X1 \cache_reg[1][1][DATA][21]  ( .D(n44), .CK(net19108), .RN(rst), .Q(
        \cache[1][1][DATA][21] ) );
  DFFR_X1 \cache_reg[1][1][DATA][20]  ( .D(n42), .CK(net19108), .RN(rst), .Q(
        \cache[1][1][DATA][20] ) );
  DFFR_X1 \cache_reg[1][1][DATA][19]  ( .D(n48), .CK(net19108), .RN(rst), .Q(
        \cache[1][1][DATA][19] ) );
  DFFR_X1 \cache_reg[1][1][DATA][18]  ( .D(n46), .CK(net19108), .RN(rst), .Q(
        \cache[1][1][DATA][18] ) );
  DFFR_X1 \cache_reg[1][1][DATA][17]  ( .D(n47), .CK(net19108), .RN(rst), .Q(
        \cache[1][1][DATA][17] ) );
  DFFR_X1 \cache_reg[1][1][DATA][16]  ( .D(n279), .CK(net19108), .RN(rst), .Q(
        \cache[1][1][DATA][16] ) );
  DFFR_X1 \cache_reg[1][1][DATA][15]  ( .D(n45), .CK(net19108), .RN(rst), .Q(
        \cache[1][1][DATA][15] ) );
  DFFR_X1 \cache_reg[1][1][DATA][14]  ( .D(n35), .CK(net19108), .RN(rst), .Q(
        \cache[1][1][DATA][14] ) );
  DFFR_X1 \cache_reg[1][1][DATA][13]  ( .D(n52), .CK(net19108), .RN(rst), .Q(
        \cache[1][1][DATA][13] ) );
  DFFR_X1 \cache_reg[1][1][DATA][12]  ( .D(n50), .CK(net19108), .RN(rst), .Q(
        \cache[1][1][DATA][12] ) );
  DFFR_X1 \cache_reg[1][1][DATA][11]  ( .D(n51), .CK(net19108), .RN(rst), .Q(
        \cache[1][1][DATA][11] ) );
  DFFR_X1 \cache_reg[1][1][DATA][10]  ( .D(n49), .CK(net19108), .RN(rst), .Q(
        \cache[1][1][DATA][10] ) );
  DFFR_X1 \cache_reg[1][1][DATA][9]  ( .D(n43), .CK(net19108), .RN(rst), .Q(
        \cache[1][1][DATA][9] ) );
  DFFR_X1 \cache_reg[1][1][DATA][8]  ( .D(n270), .CK(net19108), .RN(rst), .Q(
        \cache[1][1][DATA][8] ) );
  DFFR_X1 \cache_reg[1][1][DATA][7]  ( .D(n204), .CK(net19108), .RN(rst), .Q(
        \cache[1][1][DATA][7] ) );
  DFFR_X1 \cache_reg[1][1][DATA][6]  ( .D(n222), .CK(net19108), .RN(rst), .Q(
        \cache[1][1][DATA][6] ) );
  DFFR_X1 \cache_reg[1][1][DATA][5]  ( .D(n266), .CK(net19108), .RN(rst), .Q(
        \cache[1][1][DATA][5] ) );
  DFFR_X1 \cache_reg[1][1][DATA][4]  ( .D(n264), .CK(net19108), .RN(rst), .Q(
        \cache[1][1][DATA][4] ) );
  DFFR_X1 \cache_reg[1][1][DATA][3]  ( .D(n262), .CK(net19108), .RN(rst), .Q(
        \cache[1][1][DATA][3] ) );
  DFFR_X1 \cache_reg[1][1][DATA][2]  ( .D(n260), .CK(net19108), .RN(rst), .Q(
        \cache[1][1][DATA][2] ) );
  DFFR_X1 \cache_reg[1][1][DATA][1]  ( .D(n216), .CK(net19108), .RN(rst), .Q(
        \cache[1][1][DATA][1] ) );
  DFFR_X1 \cache_reg[1][1][DATA][0]  ( .D(n212), .CK(net19108), .RN(rst), .Q(
        \cache[1][1][DATA][0] ) );
  DFFR_X1 \cache_reg[2][1][DATA][29]  ( .D(n300), .CK(net19168), .RN(rst), .Q(
        \cache[2][1][DATA][29] ) );
  DFFR_X1 \cache_reg[2][1][DATA][28]  ( .D(n298), .CK(net19168), .RN(rst), .Q(
        \cache[2][1][DATA][28] ) );
  DFFR_X1 \cache_reg[2][1][DATA][27]  ( .D(n296), .CK(net19168), .RN(rst), .Q(
        \cache[2][1][DATA][27] ) );
  DFFR_X1 \cache_reg[2][1][DATA][26]  ( .D(n294), .CK(net19168), .RN(rst), .Q(
        \cache[2][1][DATA][26] ) );
  DFFR_X1 \cache_reg[2][1][DATA][25]  ( .D(n292), .CK(net19168), .RN(rst), .Q(
        \cache[2][1][DATA][25] ) );
  DFFR_X1 \cache_reg[2][1][DATA][24]  ( .D(n290), .CK(net19168), .RN(rst), .Q(
        \cache[2][1][DATA][24] ) );
  DFFR_X1 \cache_reg[2][1][DATA][23]  ( .D(n288), .CK(net19168), .RN(rst), .Q(
        \cache[2][1][DATA][23] ) );
  DFFR_X1 \cache_reg[2][1][DATA][22]  ( .D(n286), .CK(net19168), .RN(rst), .Q(
        \cache[2][1][DATA][22] ) );
  DFFR_X1 \cache_reg[2][1][DATA][21]  ( .D(n44), .CK(net19168), .RN(rst), .Q(
        \cache[2][1][DATA][21] ) );
  DFFR_X1 \cache_reg[2][1][DATA][20]  ( .D(n42), .CK(net19168), .RN(rst), .Q(
        \cache[2][1][DATA][20] ) );
  DFFR_X1 \cache_reg[2][1][DATA][19]  ( .D(n48), .CK(net19168), .RN(rst), .Q(
        \cache[2][1][DATA][19] ) );
  DFFR_X1 \cache_reg[2][1][DATA][18]  ( .D(n46), .CK(net19168), .RN(rst), .Q(
        \cache[2][1][DATA][18] ) );
  DFFR_X1 \cache_reg[2][1][DATA][17]  ( .D(n47), .CK(net19168), .RN(rst), .Q(
        \cache[2][1][DATA][17] ) );
  DFFR_X1 \cache_reg[2][1][DATA][16]  ( .D(n279), .CK(net19168), .RN(rst), .Q(
        \cache[2][1][DATA][16] ) );
  DFFR_X1 \cache_reg[2][1][DATA][15]  ( .D(n45), .CK(net19168), .RN(rst), .Q(
        \cache[2][1][DATA][15] ) );
  DFFR_X1 \cache_reg[2][1][DATA][14]  ( .D(n35), .CK(net19168), .RN(rst), .Q(
        \cache[2][1][DATA][14] ) );
  DFFR_X1 \cache_reg[2][1][DATA][13]  ( .D(n52), .CK(net19168), .RN(rst), .Q(
        \cache[2][1][DATA][13] ) );
  DFFR_X1 \cache_reg[2][1][DATA][12]  ( .D(n50), .CK(net19168), .RN(rst), .Q(
        \cache[2][1][DATA][12] ) );
  DFFR_X1 \cache_reg[2][1][DATA][11]  ( .D(n51), .CK(net19168), .RN(rst), .Q(
        \cache[2][1][DATA][11] ) );
  DFFR_X1 \cache_reg[2][1][DATA][10]  ( .D(n49), .CK(net19168), .RN(rst), .Q(
        \cache[2][1][DATA][10] ) );
  DFFR_X1 \cache_reg[2][1][DATA][9]  ( .D(n43), .CK(net19168), .RN(rst), .Q(
        \cache[2][1][DATA][9] ) );
  DFFR_X1 \cache_reg[2][1][DATA][8]  ( .D(n270), .CK(net19168), .RN(rst), .Q(
        \cache[2][1][DATA][8] ) );
  DFFR_X1 \cache_reg[2][1][DATA][7]  ( .D(n204), .CK(net19168), .RN(rst), .Q(
        \cache[2][1][DATA][7] ) );
  DFFR_X1 \cache_reg[2][1][DATA][6]  ( .D(n222), .CK(net19168), .RN(rst), .Q(
        \cache[2][1][DATA][6] ) );
  DFFR_X1 \cache_reg[2][1][DATA][5]  ( .D(n266), .CK(net19168), .RN(rst), .Q(
        \cache[2][1][DATA][5] ) );
  DFFR_X1 \cache_reg[2][1][DATA][4]  ( .D(n264), .CK(net19168), .RN(rst), .Q(
        \cache[2][1][DATA][4] ) );
  DFFR_X1 \cache_reg[2][1][DATA][3]  ( .D(n262), .CK(net19168), .RN(rst), .Q(
        \cache[2][1][DATA][3] ) );
  DFFR_X1 \cache_reg[2][1][DATA][2]  ( .D(n260), .CK(net19168), .RN(rst), .Q(
        \cache[2][1][DATA][2] ) );
  DFFR_X1 \cache_reg[2][1][DATA][1]  ( .D(n216), .CK(net19168), .RN(rst), .Q(
        \cache[2][1][DATA][1] ) );
  DFFR_X1 \cache_reg[2][1][DATA][0]  ( .D(n212), .CK(net19168), .RN(rst), .Q(
        \cache[2][1][DATA][0] ) );
  DFFR_X1 \cache_reg[3][1][DATA][29]  ( .D(n300), .CK(net19228), .RN(rst), .Q(
        \cache[3][1][DATA][29] ) );
  DFFR_X1 \cache_reg[3][1][DATA][28]  ( .D(n298), .CK(net19228), .RN(rst), .Q(
        \cache[3][1][DATA][28] ) );
  DFFR_X1 \cache_reg[3][1][DATA][27]  ( .D(n296), .CK(net19228), .RN(rst), .Q(
        \cache[3][1][DATA][27] ) );
  DFFR_X1 \cache_reg[3][1][DATA][26]  ( .D(n294), .CK(net19228), .RN(rst), .Q(
        \cache[3][1][DATA][26] ) );
  DFFR_X1 \cache_reg[3][1][DATA][25]  ( .D(n292), .CK(net19228), .RN(rst), .Q(
        \cache[3][1][DATA][25] ) );
  DFFR_X1 \cache_reg[3][1][DATA][24]  ( .D(n290), .CK(net19228), .RN(rst), .Q(
        \cache[3][1][DATA][24] ) );
  DFFR_X1 \cache_reg[3][1][DATA][23]  ( .D(n288), .CK(net19228), .RN(rst), .Q(
        \cache[3][1][DATA][23] ) );
  DFFR_X1 \cache_reg[3][1][DATA][22]  ( .D(n286), .CK(net19228), .RN(rst), .Q(
        \cache[3][1][DATA][22] ) );
  DFFR_X1 \cache_reg[3][1][DATA][21]  ( .D(n44), .CK(net19228), .RN(rst), .Q(
        \cache[3][1][DATA][21] ) );
  DFFR_X1 \cache_reg[3][1][DATA][20]  ( .D(n42), .CK(net19228), .RN(rst), .Q(
        \cache[3][1][DATA][20] ) );
  DFFR_X1 \cache_reg[3][1][DATA][19]  ( .D(n48), .CK(net19228), .RN(rst), .Q(
        \cache[3][1][DATA][19] ) );
  DFFR_X1 \cache_reg[3][1][DATA][18]  ( .D(n46), .CK(net19228), .RN(rst), .Q(
        \cache[3][1][DATA][18] ) );
  DFFR_X1 \cache_reg[3][1][DATA][17]  ( .D(n47), .CK(net19228), .RN(rst), .Q(
        \cache[3][1][DATA][17] ) );
  DFFR_X1 \cache_reg[3][1][DATA][16]  ( .D(n279), .CK(net19228), .RN(rst), .Q(
        \cache[3][1][DATA][16] ) );
  DFFR_X1 \cache_reg[3][1][DATA][15]  ( .D(n45), .CK(net19228), .RN(rst), .Q(
        \cache[3][1][DATA][15] ) );
  DFFR_X1 \cache_reg[3][1][DATA][14]  ( .D(n35), .CK(net19228), .RN(rst), .Q(
        \cache[3][1][DATA][14] ) );
  DFFR_X1 \cache_reg[3][1][DATA][13]  ( .D(n52), .CK(net19228), .RN(rst), .Q(
        \cache[3][1][DATA][13] ) );
  DFFR_X1 \cache_reg[3][1][DATA][12]  ( .D(n50), .CK(net19228), .RN(rst), .Q(
        \cache[3][1][DATA][12] ) );
  DFFR_X1 \cache_reg[3][1][DATA][11]  ( .D(n51), .CK(net19228), .RN(rst), .Q(
        \cache[3][1][DATA][11] ) );
  DFFR_X1 \cache_reg[3][1][DATA][10]  ( .D(n49), .CK(net19228), .RN(rst), .Q(
        \cache[3][1][DATA][10] ) );
  DFFR_X1 \cache_reg[3][1][DATA][9]  ( .D(n43), .CK(net19228), .RN(rst), .Q(
        \cache[3][1][DATA][9] ) );
  DFFR_X1 \cache_reg[3][1][DATA][8]  ( .D(n270), .CK(net19228), .RN(rst), .Q(
        \cache[3][1][DATA][8] ) );
  DFFR_X1 \cache_reg[3][1][DATA][7]  ( .D(n204), .CK(net19228), .RN(rst), .Q(
        \cache[3][1][DATA][7] ) );
  DFFR_X1 \cache_reg[3][1][DATA][6]  ( .D(n222), .CK(net19228), .RN(rst), .Q(
        \cache[3][1][DATA][6] ) );
  DFFR_X1 \cache_reg[3][1][DATA][5]  ( .D(n266), .CK(net19228), .RN(rst), .Q(
        \cache[3][1][DATA][5] ) );
  DFFR_X1 \cache_reg[3][1][DATA][4]  ( .D(n264), .CK(net19228), .RN(rst), .Q(
        \cache[3][1][DATA][4] ) );
  DFFR_X1 \cache_reg[3][1][DATA][3]  ( .D(n262), .CK(net19228), .RN(rst), .Q(
        \cache[3][1][DATA][3] ) );
  DFFR_X1 \cache_reg[3][1][DATA][2]  ( .D(n260), .CK(net19228), .RN(rst), .Q(
        \cache[3][1][DATA][2] ) );
  DFFR_X1 \cache_reg[3][1][DATA][1]  ( .D(n216), .CK(net19228), .RN(rst), .Q(
        \cache[3][1][DATA][1] ) );
  DFFR_X1 \cache_reg[3][1][DATA][0]  ( .D(n212), .CK(net19228), .RN(rst), .Q(
        \cache[3][1][DATA][0] ) );
  DFFR_X1 \cache_reg[4][1][DATA][29]  ( .D(n300), .CK(net19288), .RN(rst), .Q(
        \cache[4][1][DATA][29] ) );
  DFFR_X1 \cache_reg[4][1][DATA][28]  ( .D(n298), .CK(net19288), .RN(rst), .Q(
        \cache[4][1][DATA][28] ) );
  DFFR_X1 \cache_reg[4][1][DATA][27]  ( .D(n296), .CK(net19288), .RN(rst), .Q(
        \cache[4][1][DATA][27] ) );
  DFFR_X1 \cache_reg[4][1][DATA][26]  ( .D(n294), .CK(net19288), .RN(rst), .Q(
        \cache[4][1][DATA][26] ) );
  DFFR_X1 \cache_reg[4][1][DATA][25]  ( .D(n292), .CK(net19288), .RN(rst), .Q(
        \cache[4][1][DATA][25] ) );
  DFFR_X1 \cache_reg[4][1][DATA][24]  ( .D(n290), .CK(net19288), .RN(rst), .Q(
        \cache[4][1][DATA][24] ) );
  DFFR_X1 \cache_reg[4][1][DATA][23]  ( .D(n288), .CK(net19288), .RN(rst), .Q(
        \cache[4][1][DATA][23] ) );
  DFFR_X1 \cache_reg[4][1][DATA][22]  ( .D(n286), .CK(net19288), .RN(rst), .Q(
        \cache[4][1][DATA][22] ) );
  DFFR_X1 \cache_reg[4][1][DATA][21]  ( .D(n44), .CK(net19288), .RN(rst), .Q(
        \cache[4][1][DATA][21] ) );
  DFFR_X1 \cache_reg[4][1][DATA][20]  ( .D(n42), .CK(net19288), .RN(rst), .Q(
        \cache[4][1][DATA][20] ) );
  DFFR_X1 \cache_reg[4][1][DATA][19]  ( .D(n48), .CK(net19288), .RN(rst), .Q(
        \cache[4][1][DATA][19] ) );
  DFFR_X1 \cache_reg[4][1][DATA][18]  ( .D(n46), .CK(net19288), .RN(rst), .Q(
        \cache[4][1][DATA][18] ) );
  DFFR_X1 \cache_reg[4][1][DATA][17]  ( .D(n47), .CK(net19288), .RN(rst), .Q(
        \cache[4][1][DATA][17] ) );
  DFFR_X1 \cache_reg[4][1][DATA][16]  ( .D(n279), .CK(net19288), .RN(rst), .Q(
        \cache[4][1][DATA][16] ) );
  DFFR_X1 \cache_reg[4][1][DATA][15]  ( .D(n45), .CK(net19288), .RN(rst), .Q(
        \cache[4][1][DATA][15] ) );
  DFFR_X1 \cache_reg[4][1][DATA][14]  ( .D(n35), .CK(net19288), .RN(rst), .Q(
        \cache[4][1][DATA][14] ) );
  DFFR_X1 \cache_reg[4][1][DATA][13]  ( .D(n52), .CK(net19288), .RN(rst), .Q(
        \cache[4][1][DATA][13] ) );
  DFFR_X1 \cache_reg[4][1][DATA][12]  ( .D(n50), .CK(net19288), .RN(rst), .Q(
        \cache[4][1][DATA][12] ) );
  DFFR_X1 \cache_reg[4][1][DATA][11]  ( .D(n51), .CK(net19288), .RN(rst), .Q(
        \cache[4][1][DATA][11] ) );
  DFFR_X1 \cache_reg[4][1][DATA][10]  ( .D(n49), .CK(net19288), .RN(rst), .Q(
        \cache[4][1][DATA][10] ) );
  DFFR_X1 \cache_reg[4][1][DATA][9]  ( .D(n43), .CK(net19288), .RN(rst), .Q(
        \cache[4][1][DATA][9] ) );
  DFFR_X1 \cache_reg[4][1][DATA][8]  ( .D(n270), .CK(net19288), .RN(rst), .Q(
        \cache[4][1][DATA][8] ) );
  DFFR_X1 \cache_reg[4][1][DATA][7]  ( .D(n204), .CK(net19288), .RN(rst), .Q(
        \cache[4][1][DATA][7] ) );
  DFFR_X1 \cache_reg[4][1][DATA][6]  ( .D(n222), .CK(net19288), .RN(rst), .Q(
        \cache[4][1][DATA][6] ) );
  DFFR_X1 \cache_reg[4][1][DATA][5]  ( .D(n266), .CK(net19288), .RN(rst), .Q(
        \cache[4][1][DATA][5] ) );
  DFFR_X1 \cache_reg[4][1][DATA][4]  ( .D(n264), .CK(net19288), .RN(rst), .Q(
        \cache[4][1][DATA][4] ) );
  DFFR_X1 \cache_reg[4][1][DATA][3]  ( .D(n262), .CK(net19288), .RN(rst), .Q(
        \cache[4][1][DATA][3] ) );
  DFFR_X1 \cache_reg[4][1][DATA][2]  ( .D(n260), .CK(net19288), .RN(rst), .Q(
        \cache[4][1][DATA][2] ) );
  DFFR_X1 \cache_reg[4][1][DATA][1]  ( .D(n216), .CK(net19288), .RN(rst), .Q(
        \cache[4][1][DATA][1] ) );
  DFFR_X1 \cache_reg[4][1][DATA][0]  ( .D(n212), .CK(net19288), .RN(rst), .Q(
        \cache[4][1][DATA][0] ) );
  DFFR_X1 \cache_reg[5][1][DATA][29]  ( .D(n300), .CK(net19348), .RN(rst), .Q(
        \cache[5][1][DATA][29] ) );
  DFFR_X1 \cache_reg[5][1][DATA][28]  ( .D(n298), .CK(net19348), .RN(rst), .Q(
        \cache[5][1][DATA][28] ) );
  DFFR_X1 \cache_reg[5][1][DATA][27]  ( .D(n296), .CK(net19348), .RN(rst), .Q(
        \cache[5][1][DATA][27] ) );
  DFFR_X1 \cache_reg[5][1][DATA][26]  ( .D(n294), .CK(net19348), .RN(rst), .Q(
        \cache[5][1][DATA][26] ) );
  DFFR_X1 \cache_reg[5][1][DATA][25]  ( .D(n292), .CK(net19348), .RN(rst), .Q(
        \cache[5][1][DATA][25] ) );
  DFFR_X1 \cache_reg[5][1][DATA][24]  ( .D(n290), .CK(net19348), .RN(rst), .Q(
        \cache[5][1][DATA][24] ) );
  DFFR_X1 \cache_reg[5][1][DATA][23]  ( .D(n288), .CK(net19348), .RN(rst), .Q(
        \cache[5][1][DATA][23] ) );
  DFFR_X1 \cache_reg[5][1][DATA][22]  ( .D(n286), .CK(net19348), .RN(rst), .Q(
        \cache[5][1][DATA][22] ) );
  DFFR_X1 \cache_reg[5][1][DATA][21]  ( .D(n44), .CK(net19348), .RN(rst), .Q(
        \cache[5][1][DATA][21] ) );
  DFFR_X1 \cache_reg[5][1][DATA][20]  ( .D(n42), .CK(net19348), .RN(rst), .Q(
        \cache[5][1][DATA][20] ) );
  DFFR_X1 \cache_reg[5][1][DATA][19]  ( .D(n48), .CK(net19348), .RN(rst), .Q(
        \cache[5][1][DATA][19] ) );
  DFFR_X1 \cache_reg[5][1][DATA][18]  ( .D(n46), .CK(net19348), .RN(rst), .Q(
        \cache[5][1][DATA][18] ) );
  DFFR_X1 \cache_reg[5][1][DATA][17]  ( .D(n47), .CK(net19348), .RN(rst), .Q(
        \cache[5][1][DATA][17] ) );
  DFFR_X1 \cache_reg[5][1][DATA][16]  ( .D(n279), .CK(net19348), .RN(rst), .Q(
        \cache[5][1][DATA][16] ) );
  DFFR_X1 \cache_reg[5][1][DATA][15]  ( .D(n45), .CK(net19348), .RN(rst), .Q(
        \cache[5][1][DATA][15] ) );
  DFFR_X1 \cache_reg[5][1][DATA][14]  ( .D(n35), .CK(net19348), .RN(rst), .Q(
        \cache[5][1][DATA][14] ) );
  DFFR_X1 \cache_reg[5][1][DATA][13]  ( .D(n52), .CK(net19348), .RN(rst), .Q(
        \cache[5][1][DATA][13] ) );
  DFFR_X1 \cache_reg[5][1][DATA][12]  ( .D(n50), .CK(net19348), .RN(rst), .Q(
        \cache[5][1][DATA][12] ) );
  DFFR_X1 \cache_reg[5][1][DATA][11]  ( .D(n51), .CK(net19348), .RN(rst), .Q(
        \cache[5][1][DATA][11] ) );
  DFFR_X1 \cache_reg[5][1][DATA][10]  ( .D(n49), .CK(net19348), .RN(rst), .Q(
        \cache[5][1][DATA][10] ) );
  DFFR_X1 \cache_reg[5][1][DATA][9]  ( .D(n43), .CK(net19348), .RN(rst), .Q(
        \cache[5][1][DATA][9] ) );
  DFFR_X1 \cache_reg[5][1][DATA][8]  ( .D(n270), .CK(net19348), .RN(rst), .Q(
        \cache[5][1][DATA][8] ) );
  DFFR_X1 \cache_reg[5][1][DATA][7]  ( .D(n204), .CK(net19348), .RN(rst), .Q(
        \cache[5][1][DATA][7] ) );
  DFFR_X1 \cache_reg[5][1][DATA][6]  ( .D(n222), .CK(net19348), .RN(rst), .Q(
        \cache[5][1][DATA][6] ) );
  DFFR_X1 \cache_reg[5][1][DATA][5]  ( .D(n266), .CK(net19348), .RN(rst), .Q(
        \cache[5][1][DATA][5] ) );
  DFFR_X1 \cache_reg[5][1][DATA][4]  ( .D(n264), .CK(net19348), .RN(rst), .Q(
        \cache[5][1][DATA][4] ) );
  DFFR_X1 \cache_reg[5][1][DATA][3]  ( .D(n262), .CK(net19348), .RN(rst), .Q(
        \cache[5][1][DATA][3] ) );
  DFFR_X1 \cache_reg[5][1][DATA][2]  ( .D(n260), .CK(net19348), .RN(rst), .Q(
        \cache[5][1][DATA][2] ) );
  DFFR_X1 \cache_reg[5][1][DATA][1]  ( .D(n216), .CK(net19348), .RN(rst), .Q(
        \cache[5][1][DATA][1] ) );
  DFFR_X1 \cache_reg[5][1][DATA][0]  ( .D(n212), .CK(net19348), .RN(rst), .Q(
        \cache[5][1][DATA][0] ) );
  DFFR_X1 \cache_reg[6][1][DATA][29]  ( .D(n300), .CK(net19408), .RN(rst), .Q(
        \cache[6][1][DATA][29] ) );
  DFFR_X1 \cache_reg[6][1][DATA][28]  ( .D(n298), .CK(net19408), .RN(rst), .Q(
        \cache[6][1][DATA][28] ) );
  DFFR_X1 \cache_reg[6][1][DATA][27]  ( .D(n296), .CK(net19408), .RN(rst), .Q(
        \cache[6][1][DATA][27] ) );
  DFFR_X1 \cache_reg[6][1][DATA][26]  ( .D(n294), .CK(net19408), .RN(rst), .Q(
        \cache[6][1][DATA][26] ) );
  DFFR_X1 \cache_reg[6][1][DATA][25]  ( .D(n292), .CK(net19408), .RN(rst), .Q(
        \cache[6][1][DATA][25] ) );
  DFFR_X1 \cache_reg[6][1][DATA][24]  ( .D(n290), .CK(net19408), .RN(rst), .Q(
        \cache[6][1][DATA][24] ) );
  DFFR_X1 \cache_reg[6][1][DATA][23]  ( .D(n288), .CK(net19408), .RN(rst), .Q(
        \cache[6][1][DATA][23] ) );
  DFFR_X1 \cache_reg[6][1][DATA][22]  ( .D(n286), .CK(net19408), .RN(rst), .Q(
        \cache[6][1][DATA][22] ) );
  DFFR_X1 \cache_reg[6][1][DATA][21]  ( .D(n44), .CK(net19408), .RN(rst), .Q(
        \cache[6][1][DATA][21] ) );
  DFFR_X1 \cache_reg[6][1][DATA][20]  ( .D(n42), .CK(net19408), .RN(rst), .Q(
        \cache[6][1][DATA][20] ) );
  DFFR_X1 \cache_reg[6][1][DATA][19]  ( .D(n48), .CK(net19408), .RN(rst), .Q(
        \cache[6][1][DATA][19] ) );
  DFFR_X1 \cache_reg[6][1][DATA][18]  ( .D(n46), .CK(net19408), .RN(rst), .Q(
        \cache[6][1][DATA][18] ) );
  DFFR_X1 \cache_reg[6][1][DATA][17]  ( .D(n47), .CK(net19408), .RN(rst), .Q(
        \cache[6][1][DATA][17] ) );
  DFFR_X1 \cache_reg[6][1][DATA][16]  ( .D(n279), .CK(net19408), .RN(rst), .Q(
        \cache[6][1][DATA][16] ) );
  DFFR_X1 \cache_reg[6][1][DATA][15]  ( .D(n45), .CK(net19408), .RN(rst), .Q(
        \cache[6][1][DATA][15] ) );
  DFFR_X1 \cache_reg[6][1][DATA][14]  ( .D(n35), .CK(net19408), .RN(rst), .Q(
        \cache[6][1][DATA][14] ) );
  DFFR_X1 \cache_reg[6][1][DATA][13]  ( .D(n52), .CK(net19408), .RN(rst), .Q(
        \cache[6][1][DATA][13] ) );
  DFFR_X1 \cache_reg[6][1][DATA][12]  ( .D(n50), .CK(net19408), .RN(rst), .Q(
        \cache[6][1][DATA][12] ) );
  DFFR_X1 \cache_reg[6][1][DATA][11]  ( .D(n51), .CK(net19408), .RN(rst), .Q(
        \cache[6][1][DATA][11] ) );
  DFFR_X1 \cache_reg[6][1][DATA][10]  ( .D(n49), .CK(net19408), .RN(rst), .Q(
        \cache[6][1][DATA][10] ) );
  DFFR_X1 \cache_reg[6][1][DATA][9]  ( .D(n43), .CK(net19408), .RN(rst), .Q(
        \cache[6][1][DATA][9] ) );
  DFFR_X1 \cache_reg[6][1][DATA][8]  ( .D(n270), .CK(net19408), .RN(rst), .Q(
        \cache[6][1][DATA][8] ) );
  DFFR_X1 \cache_reg[6][1][DATA][7]  ( .D(n204), .CK(net19408), .RN(rst), .Q(
        \cache[6][1][DATA][7] ) );
  DFFR_X1 \cache_reg[6][1][DATA][6]  ( .D(n222), .CK(net19408), .RN(rst), .Q(
        \cache[6][1][DATA][6] ) );
  DFFR_X1 \cache_reg[6][1][DATA][5]  ( .D(n266), .CK(net19408), .RN(rst), .Q(
        \cache[6][1][DATA][5] ) );
  DFFR_X1 \cache_reg[6][1][DATA][4]  ( .D(n264), .CK(net19408), .RN(rst), .Q(
        \cache[6][1][DATA][4] ) );
  DFFR_X1 \cache_reg[6][1][DATA][3]  ( .D(n262), .CK(net19408), .RN(rst), .Q(
        \cache[6][1][DATA][3] ) );
  DFFR_X1 \cache_reg[6][1][DATA][2]  ( .D(n260), .CK(net19408), .RN(rst), .Q(
        \cache[6][1][DATA][2] ) );
  DFFR_X1 \cache_reg[6][1][DATA][1]  ( .D(n216), .CK(net19408), .RN(rst), .Q(
        \cache[6][1][DATA][1] ) );
  DFFR_X1 \cache_reg[6][1][DATA][0]  ( .D(n212), .CK(net19408), .RN(rst), .Q(
        \cache[6][1][DATA][0] ) );
  DFFR_X1 \cache_reg[7][1][DATA][29]  ( .D(n300), .CK(net19468), .RN(rst), .Q(
        \cache[7][1][DATA][29] ) );
  DFFR_X1 \cache_reg[7][1][DATA][28]  ( .D(n298), .CK(net19468), .RN(rst), .Q(
        \cache[7][1][DATA][28] ) );
  DFFR_X1 \cache_reg[7][1][DATA][27]  ( .D(n296), .CK(net19468), .RN(rst), .Q(
        \cache[7][1][DATA][27] ) );
  DFFR_X1 \cache_reg[7][1][DATA][26]  ( .D(n294), .CK(net19468), .RN(rst), .Q(
        \cache[7][1][DATA][26] ) );
  DFFR_X1 \cache_reg[7][1][DATA][25]  ( .D(n292), .CK(net19468), .RN(rst), .Q(
        \cache[7][1][DATA][25] ) );
  DFFR_X1 \cache_reg[7][1][DATA][24]  ( .D(n290), .CK(net19468), .RN(rst), .Q(
        \cache[7][1][DATA][24] ) );
  DFFR_X1 \cache_reg[7][1][DATA][23]  ( .D(n288), .CK(net19468), .RN(rst), .Q(
        \cache[7][1][DATA][23] ) );
  DFFR_X1 \cache_reg[7][1][DATA][22]  ( .D(n286), .CK(net19468), .RN(rst), .Q(
        \cache[7][1][DATA][22] ) );
  DFFR_X1 \cache_reg[7][1][DATA][21]  ( .D(n44), .CK(net19468), .RN(rst), .Q(
        \cache[7][1][DATA][21] ) );
  DFFR_X1 \cache_reg[7][1][DATA][20]  ( .D(n42), .CK(net19468), .RN(rst), .Q(
        \cache[7][1][DATA][20] ) );
  DFFR_X1 \cache_reg[7][1][DATA][19]  ( .D(n48), .CK(net19468), .RN(rst), .Q(
        \cache[7][1][DATA][19] ) );
  DFFR_X1 \cache_reg[7][1][DATA][18]  ( .D(n46), .CK(net19468), .RN(rst), .Q(
        \cache[7][1][DATA][18] ) );
  DFFR_X1 \cache_reg[7][1][DATA][17]  ( .D(n47), .CK(net19468), .RN(rst), .Q(
        \cache[7][1][DATA][17] ) );
  DFFR_X1 \cache_reg[7][1][DATA][16]  ( .D(n279), .CK(net19468), .RN(rst), .Q(
        \cache[7][1][DATA][16] ) );
  DFFR_X1 \cache_reg[7][1][DATA][15]  ( .D(n45), .CK(net19468), .RN(rst), .Q(
        \cache[7][1][DATA][15] ) );
  DFFR_X1 \cache_reg[7][1][DATA][14]  ( .D(n35), .CK(net19468), .RN(rst), .Q(
        \cache[7][1][DATA][14] ) );
  DFFR_X1 \cache_reg[7][1][DATA][13]  ( .D(n52), .CK(net19468), .RN(rst), .Q(
        \cache[7][1][DATA][13] ) );
  DFFR_X1 \cache_reg[7][1][DATA][12]  ( .D(n50), .CK(net19468), .RN(rst), .Q(
        \cache[7][1][DATA][12] ) );
  DFFR_X1 \cache_reg[7][1][DATA][11]  ( .D(n51), .CK(net19468), .RN(rst), .Q(
        \cache[7][1][DATA][11] ) );
  DFFR_X1 \cache_reg[7][1][DATA][10]  ( .D(n49), .CK(net19468), .RN(rst), .Q(
        \cache[7][1][DATA][10] ) );
  DFFR_X1 \cache_reg[7][1][DATA][9]  ( .D(n43), .CK(net19468), .RN(rst), .Q(
        \cache[7][1][DATA][9] ) );
  DFFR_X1 \cache_reg[7][1][DATA][8]  ( .D(n270), .CK(net19468), .RN(rst), .Q(
        \cache[7][1][DATA][8] ) );
  DFFR_X1 \cache_reg[7][1][DATA][7]  ( .D(n204), .CK(net19468), .RN(rst), .Q(
        \cache[7][1][DATA][7] ) );
  DFFR_X1 \cache_reg[7][1][DATA][6]  ( .D(n222), .CK(net19468), .RN(rst), .Q(
        \cache[7][1][DATA][6] ) );
  DFFR_X1 \cache_reg[7][1][DATA][5]  ( .D(n266), .CK(net19468), .RN(rst), .Q(
        \cache[7][1][DATA][5] ) );
  DFFR_X1 \cache_reg[7][1][DATA][4]  ( .D(n264), .CK(net19468), .RN(rst), .Q(
        \cache[7][1][DATA][4] ) );
  DFFR_X1 \cache_reg[7][1][DATA][3]  ( .D(n262), .CK(net19468), .RN(rst), .Q(
        \cache[7][1][DATA][3] ) );
  DFFR_X1 \cache_reg[7][1][DATA][2]  ( .D(n260), .CK(net19468), .RN(rst), .Q(
        \cache[7][1][DATA][2] ) );
  DFFR_X1 \cache_reg[7][1][DATA][1]  ( .D(n216), .CK(net19468), .RN(rst), .Q(
        \cache[7][1][DATA][1] ) );
  DFFR_X1 \cache_reg[7][1][DATA][0]  ( .D(n212), .CK(net19468), .RN(rst), .Q(
        \cache[7][1][DATA][0] ) );
  DFFR_X1 \cache_reg[0][2][DATA][29]  ( .D(n300), .CK(net19063), .RN(rst), .Q(
        \cache[0][2][DATA][29] ) );
  DFFR_X1 \cache_reg[0][2][DATA][28]  ( .D(n298), .CK(net19063), .RN(rst), .Q(
        \cache[0][2][DATA][28] ) );
  DFFR_X1 \cache_reg[0][2][DATA][27]  ( .D(n296), .CK(net19063), .RN(rst), .Q(
        \cache[0][2][DATA][27] ) );
  DFFR_X1 \cache_reg[0][2][DATA][26]  ( .D(n294), .CK(net19063), .RN(rst), .Q(
        \cache[0][2][DATA][26] ) );
  DFFR_X1 \cache_reg[0][2][DATA][25]  ( .D(n292), .CK(net19063), .RN(rst), .Q(
        \cache[0][2][DATA][25] ) );
  DFFR_X1 \cache_reg[0][2][DATA][24]  ( .D(n290), .CK(net19063), .RN(rst), .Q(
        \cache[0][2][DATA][24] ) );
  DFFR_X1 \cache_reg[0][2][DATA][23]  ( .D(n288), .CK(net19063), .RN(rst), .Q(
        \cache[0][2][DATA][23] ) );
  DFFR_X1 \cache_reg[0][2][DATA][22]  ( .D(n286), .CK(net19063), .RN(rst), .Q(
        \cache[0][2][DATA][22] ) );
  DFFR_X1 \cache_reg[0][2][DATA][21]  ( .D(n44), .CK(net19063), .RN(rst), .Q(
        \cache[0][2][DATA][21] ) );
  DFFR_X1 \cache_reg[0][2][DATA][20]  ( .D(n42), .CK(net19063), .RN(rst), .Q(
        \cache[0][2][DATA][20] ) );
  DFFR_X1 \cache_reg[0][2][DATA][19]  ( .D(n48), .CK(net19063), .RN(rst), .Q(
        \cache[0][2][DATA][19] ) );
  DFFR_X1 \cache_reg[0][2][DATA][18]  ( .D(n46), .CK(net19063), .RN(rst), .Q(
        \cache[0][2][DATA][18] ) );
  DFFR_X1 \cache_reg[0][2][DATA][17]  ( .D(n47), .CK(net19063), .RN(rst), .Q(
        \cache[0][2][DATA][17] ) );
  DFFR_X1 \cache_reg[0][2][DATA][16]  ( .D(n279), .CK(net19063), .RN(rst), .Q(
        \cache[0][2][DATA][16] ) );
  DFFR_X1 \cache_reg[0][2][DATA][15]  ( .D(n45), .CK(net19063), .RN(rst), .Q(
        \cache[0][2][DATA][15] ) );
  DFFR_X1 \cache_reg[0][2][DATA][14]  ( .D(n35), .CK(net19063), .RN(rst), .Q(
        \cache[0][2][DATA][14] ) );
  DFFR_X1 \cache_reg[0][2][DATA][13]  ( .D(n52), .CK(net19063), .RN(rst), .Q(
        \cache[0][2][DATA][13] ) );
  DFFR_X1 \cache_reg[0][2][DATA][12]  ( .D(n50), .CK(net19063), .RN(rst), .Q(
        \cache[0][2][DATA][12] ) );
  DFFR_X1 \cache_reg[0][2][DATA][11]  ( .D(n51), .CK(net19063), .RN(rst), .Q(
        \cache[0][2][DATA][11] ) );
  DFFR_X1 \cache_reg[0][2][DATA][10]  ( .D(n49), .CK(net19063), .RN(rst), .Q(
        \cache[0][2][DATA][10] ) );
  DFFR_X1 \cache_reg[0][2][DATA][9]  ( .D(n43), .CK(net19063), .RN(rst), .Q(
        \cache[0][2][DATA][9] ) );
  DFFR_X1 \cache_reg[0][2][DATA][8]  ( .D(n270), .CK(net19063), .RN(rst), .Q(
        \cache[0][2][DATA][8] ) );
  DFFR_X1 \cache_reg[0][2][DATA][7]  ( .D(n204), .CK(net19063), .RN(rst), .Q(
        \cache[0][2][DATA][7] ) );
  DFFR_X1 \cache_reg[0][2][DATA][6]  ( .D(n222), .CK(net19063), .RN(rst), .Q(
        \cache[0][2][DATA][6] ) );
  DFFR_X1 \cache_reg[0][2][DATA][5]  ( .D(n266), .CK(net19063), .RN(rst), .Q(
        \cache[0][2][DATA][5] ) );
  DFFR_X1 \cache_reg[0][2][DATA][4]  ( .D(n264), .CK(net19063), .RN(rst), .Q(
        \cache[0][2][DATA][4] ) );
  DFFR_X1 \cache_reg[0][2][DATA][3]  ( .D(n262), .CK(net19063), .RN(rst), .Q(
        \cache[0][2][DATA][3] ) );
  DFFR_X1 \cache_reg[0][2][DATA][2]  ( .D(n260), .CK(net19063), .RN(rst), .Q(
        \cache[0][2][DATA][2] ) );
  DFFR_X1 \cache_reg[0][2][DATA][1]  ( .D(n216), .CK(net19063), .RN(rst), .Q(
        \cache[0][2][DATA][1] ) );
  DFFR_X1 \cache_reg[0][2][DATA][0]  ( .D(n212), .CK(net19063), .RN(rst), .Q(
        \cache[0][2][DATA][0] ) );
  DFFR_X1 \cache_reg[1][2][DATA][29]  ( .D(n300), .CK(net19123), .RN(rst), .Q(
        \cache[1][2][DATA][29] ) );
  DFFR_X1 \cache_reg[1][2][DATA][28]  ( .D(n298), .CK(net19123), .RN(rst), .Q(
        \cache[1][2][DATA][28] ) );
  DFFR_X1 \cache_reg[1][2][DATA][27]  ( .D(n296), .CK(net19123), .RN(rst), .Q(
        \cache[1][2][DATA][27] ) );
  DFFR_X1 \cache_reg[1][2][DATA][26]  ( .D(n294), .CK(net19123), .RN(rst), .Q(
        \cache[1][2][DATA][26] ) );
  DFFR_X1 \cache_reg[1][2][DATA][25]  ( .D(n292), .CK(net19123), .RN(rst), .Q(
        \cache[1][2][DATA][25] ) );
  DFFR_X1 \cache_reg[1][2][DATA][24]  ( .D(n290), .CK(net19123), .RN(rst), .Q(
        \cache[1][2][DATA][24] ) );
  DFFR_X1 \cache_reg[1][2][DATA][23]  ( .D(n288), .CK(net19123), .RN(rst), .Q(
        \cache[1][2][DATA][23] ) );
  DFFR_X1 \cache_reg[1][2][DATA][22]  ( .D(n286), .CK(net19123), .RN(rst), .Q(
        \cache[1][2][DATA][22] ) );
  DFFR_X1 \cache_reg[1][2][DATA][21]  ( .D(n44), .CK(net19123), .RN(rst), .Q(
        \cache[1][2][DATA][21] ) );
  DFFR_X1 \cache_reg[1][2][DATA][20]  ( .D(n42), .CK(net19123), .RN(rst), .Q(
        \cache[1][2][DATA][20] ) );
  DFFR_X1 \cache_reg[1][2][DATA][19]  ( .D(n48), .CK(net19123), .RN(rst), .Q(
        \cache[1][2][DATA][19] ) );
  DFFR_X1 \cache_reg[1][2][DATA][18]  ( .D(n46), .CK(net19123), .RN(rst), .Q(
        \cache[1][2][DATA][18] ) );
  DFFR_X1 \cache_reg[1][2][DATA][17]  ( .D(n47), .CK(net19123), .RN(rst), .Q(
        \cache[1][2][DATA][17] ) );
  DFFR_X1 \cache_reg[1][2][DATA][16]  ( .D(n279), .CK(net19123), .RN(rst), .Q(
        \cache[1][2][DATA][16] ) );
  DFFR_X1 \cache_reg[1][2][DATA][15]  ( .D(n45), .CK(net19123), .RN(rst), .Q(
        \cache[1][2][DATA][15] ) );
  DFFR_X1 \cache_reg[1][2][DATA][14]  ( .D(n35), .CK(net19123), .RN(rst), .Q(
        \cache[1][2][DATA][14] ) );
  DFFR_X1 \cache_reg[1][2][DATA][13]  ( .D(n52), .CK(net19123), .RN(rst), .Q(
        \cache[1][2][DATA][13] ) );
  DFFR_X1 \cache_reg[1][2][DATA][12]  ( .D(n50), .CK(net19123), .RN(rst), .Q(
        \cache[1][2][DATA][12] ) );
  DFFR_X1 \cache_reg[1][2][DATA][11]  ( .D(n51), .CK(net19123), .RN(rst), .Q(
        \cache[1][2][DATA][11] ) );
  DFFR_X1 \cache_reg[1][2][DATA][10]  ( .D(n49), .CK(net19123), .RN(rst), .Q(
        \cache[1][2][DATA][10] ) );
  DFFR_X1 \cache_reg[1][2][DATA][9]  ( .D(n43), .CK(net19123), .RN(rst), .Q(
        \cache[1][2][DATA][9] ) );
  DFFR_X1 \cache_reg[1][2][DATA][8]  ( .D(n270), .CK(net19123), .RN(rst), .Q(
        \cache[1][2][DATA][8] ) );
  DFFR_X1 \cache_reg[1][2][DATA][7]  ( .D(n204), .CK(net19123), .RN(rst), .Q(
        \cache[1][2][DATA][7] ) );
  DFFR_X1 \cache_reg[1][2][DATA][6]  ( .D(n222), .CK(net19123), .RN(rst), .Q(
        \cache[1][2][DATA][6] ) );
  DFFR_X1 \cache_reg[1][2][DATA][5]  ( .D(n266), .CK(net19123), .RN(rst), .Q(
        \cache[1][2][DATA][5] ) );
  DFFR_X1 \cache_reg[1][2][DATA][4]  ( .D(n264), .CK(net19123), .RN(rst), .Q(
        \cache[1][2][DATA][4] ) );
  DFFR_X1 \cache_reg[1][2][DATA][3]  ( .D(n262), .CK(net19123), .RN(rst), .Q(
        \cache[1][2][DATA][3] ) );
  DFFR_X1 \cache_reg[1][2][DATA][2]  ( .D(n260), .CK(net19123), .RN(rst), .Q(
        \cache[1][2][DATA][2] ) );
  DFFR_X1 \cache_reg[1][2][DATA][1]  ( .D(n216), .CK(net19123), .RN(rst), .Q(
        \cache[1][2][DATA][1] ) );
  DFFR_X1 \cache_reg[1][2][DATA][0]  ( .D(n212), .CK(net19123), .RN(rst), .Q(
        \cache[1][2][DATA][0] ) );
  DFFR_X1 \cache_reg[2][2][DATA][29]  ( .D(n300), .CK(net19183), .RN(rst), .Q(
        \cache[2][2][DATA][29] ) );
  DFFR_X1 \cache_reg[2][2][DATA][28]  ( .D(n298), .CK(net19183), .RN(rst), .Q(
        \cache[2][2][DATA][28] ) );
  DFFR_X1 \cache_reg[2][2][DATA][27]  ( .D(n296), .CK(net19183), .RN(rst), .Q(
        \cache[2][2][DATA][27] ) );
  DFFR_X1 \cache_reg[2][2][DATA][26]  ( .D(n294), .CK(net19183), .RN(rst), .Q(
        \cache[2][2][DATA][26] ) );
  DFFR_X1 \cache_reg[2][2][DATA][25]  ( .D(n292), .CK(net19183), .RN(rst), .Q(
        \cache[2][2][DATA][25] ) );
  DFFR_X1 \cache_reg[2][2][DATA][24]  ( .D(n290), .CK(net19183), .RN(rst), .Q(
        \cache[2][2][DATA][24] ) );
  DFFR_X1 \cache_reg[2][2][DATA][23]  ( .D(n288), .CK(net19183), .RN(rst), .Q(
        \cache[2][2][DATA][23] ) );
  DFFR_X1 \cache_reg[2][2][DATA][22]  ( .D(n286), .CK(net19183), .RN(rst), .Q(
        \cache[2][2][DATA][22] ) );
  DFFR_X1 \cache_reg[2][2][DATA][21]  ( .D(n44), .CK(net19183), .RN(rst), .Q(
        \cache[2][2][DATA][21] ) );
  DFFR_X1 \cache_reg[2][2][DATA][20]  ( .D(n42), .CK(net19183), .RN(rst), .Q(
        \cache[2][2][DATA][20] ) );
  DFFR_X1 \cache_reg[2][2][DATA][19]  ( .D(n48), .CK(net19183), .RN(rst), .Q(
        \cache[2][2][DATA][19] ) );
  DFFR_X1 \cache_reg[2][2][DATA][18]  ( .D(n46), .CK(net19183), .RN(rst), .Q(
        \cache[2][2][DATA][18] ) );
  DFFR_X1 \cache_reg[2][2][DATA][17]  ( .D(n47), .CK(net19183), .RN(rst), .Q(
        \cache[2][2][DATA][17] ) );
  DFFR_X1 \cache_reg[2][2][DATA][16]  ( .D(n279), .CK(net19183), .RN(rst), .Q(
        \cache[2][2][DATA][16] ) );
  DFFR_X1 \cache_reg[2][2][DATA][15]  ( .D(n45), .CK(net19183), .RN(rst), .Q(
        \cache[2][2][DATA][15] ) );
  DFFR_X1 \cache_reg[2][2][DATA][14]  ( .D(n35), .CK(net19183), .RN(rst), .Q(
        \cache[2][2][DATA][14] ) );
  DFFR_X1 \cache_reg[2][2][DATA][13]  ( .D(n52), .CK(net19183), .RN(rst), .Q(
        \cache[2][2][DATA][13] ) );
  DFFR_X1 \cache_reg[2][2][DATA][12]  ( .D(n50), .CK(net19183), .RN(rst), .Q(
        \cache[2][2][DATA][12] ) );
  DFFR_X1 \cache_reg[2][2][DATA][11]  ( .D(n51), .CK(net19183), .RN(rst), .Q(
        \cache[2][2][DATA][11] ) );
  DFFR_X1 \cache_reg[2][2][DATA][10]  ( .D(n49), .CK(net19183), .RN(rst), .Q(
        \cache[2][2][DATA][10] ) );
  DFFR_X1 \cache_reg[2][2][DATA][9]  ( .D(n43), .CK(net19183), .RN(rst), .Q(
        \cache[2][2][DATA][9] ) );
  DFFR_X1 \cache_reg[2][2][DATA][8]  ( .D(n270), .CK(net19183), .RN(rst), .Q(
        \cache[2][2][DATA][8] ) );
  DFFR_X1 \cache_reg[2][2][DATA][7]  ( .D(n204), .CK(net19183), .RN(rst), .Q(
        \cache[2][2][DATA][7] ) );
  DFFR_X1 \cache_reg[2][2][DATA][6]  ( .D(n222), .CK(net19183), .RN(rst), .Q(
        \cache[2][2][DATA][6] ) );
  DFFR_X1 \cache_reg[2][2][DATA][5]  ( .D(n266), .CK(net19183), .RN(rst), .Q(
        \cache[2][2][DATA][5] ) );
  DFFR_X1 \cache_reg[2][2][DATA][4]  ( .D(n264), .CK(net19183), .RN(rst), .Q(
        \cache[2][2][DATA][4] ) );
  DFFR_X1 \cache_reg[2][2][DATA][3]  ( .D(n262), .CK(net19183), .RN(rst), .Q(
        \cache[2][2][DATA][3] ) );
  DFFR_X1 \cache_reg[2][2][DATA][2]  ( .D(n260), .CK(net19183), .RN(rst), .Q(
        \cache[2][2][DATA][2] ) );
  DFFR_X1 \cache_reg[2][2][DATA][1]  ( .D(n216), .CK(net19183), .RN(rst), .Q(
        \cache[2][2][DATA][1] ) );
  DFFR_X1 \cache_reg[2][2][DATA][0]  ( .D(n212), .CK(net19183), .RN(rst), .Q(
        \cache[2][2][DATA][0] ) );
  DFFR_X1 \cache_reg[3][2][DATA][29]  ( .D(n300), .CK(net19243), .RN(rst), .Q(
        \cache[3][2][DATA][29] ) );
  DFFR_X1 \cache_reg[3][2][DATA][28]  ( .D(n298), .CK(net19243), .RN(rst), .Q(
        \cache[3][2][DATA][28] ) );
  DFFR_X1 \cache_reg[3][2][DATA][27]  ( .D(n296), .CK(net19243), .RN(rst), .Q(
        \cache[3][2][DATA][27] ) );
  DFFR_X1 \cache_reg[3][2][DATA][26]  ( .D(n294), .CK(net19243), .RN(rst), .Q(
        \cache[3][2][DATA][26] ) );
  DFFR_X1 \cache_reg[3][2][DATA][25]  ( .D(n292), .CK(net19243), .RN(rst), .Q(
        \cache[3][2][DATA][25] ) );
  DFFR_X1 \cache_reg[3][2][DATA][24]  ( .D(n290), .CK(net19243), .RN(rst), .Q(
        \cache[3][2][DATA][24] ) );
  DFFR_X1 \cache_reg[3][2][DATA][23]  ( .D(n288), .CK(net19243), .RN(rst), .Q(
        \cache[3][2][DATA][23] ) );
  DFFR_X1 \cache_reg[3][2][DATA][22]  ( .D(n286), .CK(net19243), .RN(rst), .Q(
        \cache[3][2][DATA][22] ) );
  DFFR_X1 \cache_reg[3][2][DATA][21]  ( .D(n44), .CK(net19243), .RN(rst), .Q(
        \cache[3][2][DATA][21] ) );
  DFFR_X1 \cache_reg[3][2][DATA][20]  ( .D(n42), .CK(net19243), .RN(rst), .Q(
        \cache[3][2][DATA][20] ) );
  DFFR_X1 \cache_reg[3][2][DATA][19]  ( .D(n48), .CK(net19243), .RN(rst), .Q(
        \cache[3][2][DATA][19] ) );
  DFFR_X1 \cache_reg[3][2][DATA][18]  ( .D(n46), .CK(net19243), .RN(rst), .Q(
        \cache[3][2][DATA][18] ) );
  DFFR_X1 \cache_reg[3][2][DATA][17]  ( .D(n47), .CK(net19243), .RN(rst), .Q(
        \cache[3][2][DATA][17] ) );
  DFFR_X1 \cache_reg[3][2][DATA][16]  ( .D(n279), .CK(net19243), .RN(rst), .Q(
        \cache[3][2][DATA][16] ) );
  DFFR_X1 \cache_reg[3][2][DATA][15]  ( .D(n45), .CK(net19243), .RN(rst), .Q(
        \cache[3][2][DATA][15] ) );
  DFFR_X1 \cache_reg[3][2][DATA][14]  ( .D(n35), .CK(net19243), .RN(rst), .Q(
        \cache[3][2][DATA][14] ) );
  DFFR_X1 \cache_reg[3][2][DATA][13]  ( .D(n52), .CK(net19243), .RN(rst), .Q(
        \cache[3][2][DATA][13] ) );
  DFFR_X1 \cache_reg[3][2][DATA][12]  ( .D(n50), .CK(net19243), .RN(rst), .Q(
        \cache[3][2][DATA][12] ) );
  DFFR_X1 \cache_reg[3][2][DATA][11]  ( .D(n51), .CK(net19243), .RN(rst), .Q(
        \cache[3][2][DATA][11] ) );
  DFFR_X1 \cache_reg[3][2][DATA][10]  ( .D(n49), .CK(net19243), .RN(rst), .Q(
        \cache[3][2][DATA][10] ) );
  DFFR_X1 \cache_reg[3][2][DATA][9]  ( .D(n43), .CK(net19243), .RN(rst), .Q(
        \cache[3][2][DATA][9] ) );
  DFFR_X1 \cache_reg[3][2][DATA][8]  ( .D(n270), .CK(net19243), .RN(rst), .Q(
        \cache[3][2][DATA][8] ) );
  DFFR_X1 \cache_reg[3][2][DATA][7]  ( .D(n204), .CK(net19243), .RN(rst), .Q(
        \cache[3][2][DATA][7] ) );
  DFFR_X1 \cache_reg[3][2][DATA][6]  ( .D(n222), .CK(net19243), .RN(rst), .Q(
        \cache[3][2][DATA][6] ) );
  DFFR_X1 \cache_reg[3][2][DATA][5]  ( .D(n266), .CK(net19243), .RN(rst), .Q(
        \cache[3][2][DATA][5] ) );
  DFFR_X1 \cache_reg[3][2][DATA][4]  ( .D(n264), .CK(net19243), .RN(rst), .Q(
        \cache[3][2][DATA][4] ) );
  DFFR_X1 \cache_reg[3][2][DATA][3]  ( .D(n262), .CK(net19243), .RN(rst), .Q(
        \cache[3][2][DATA][3] ) );
  DFFR_X1 \cache_reg[3][2][DATA][2]  ( .D(n260), .CK(net19243), .RN(rst), .Q(
        \cache[3][2][DATA][2] ) );
  DFFR_X1 \cache_reg[3][2][DATA][1]  ( .D(n216), .CK(net19243), .RN(rst), .Q(
        \cache[3][2][DATA][1] ) );
  DFFR_X1 \cache_reg[3][2][DATA][0]  ( .D(n212), .CK(net19243), .RN(rst), .Q(
        \cache[3][2][DATA][0] ) );
  DFFR_X1 \cache_reg[4][2][DATA][29]  ( .D(n300), .CK(net19303), .RN(rst), .Q(
        \cache[4][2][DATA][29] ) );
  DFFR_X1 \cache_reg[4][2][DATA][28]  ( .D(n298), .CK(net19303), .RN(rst), .Q(
        \cache[4][2][DATA][28] ) );
  DFFR_X1 \cache_reg[4][2][DATA][27]  ( .D(n296), .CK(net19303), .RN(rst), .Q(
        \cache[4][2][DATA][27] ) );
  DFFR_X1 \cache_reg[4][2][DATA][26]  ( .D(n294), .CK(net19303), .RN(rst), .Q(
        \cache[4][2][DATA][26] ) );
  DFFR_X1 \cache_reg[4][2][DATA][25]  ( .D(n292), .CK(net19303), .RN(rst), .Q(
        \cache[4][2][DATA][25] ) );
  DFFR_X1 \cache_reg[4][2][DATA][24]  ( .D(n290), .CK(net19303), .RN(rst), .Q(
        \cache[4][2][DATA][24] ) );
  DFFR_X1 \cache_reg[4][2][DATA][23]  ( .D(n288), .CK(net19303), .RN(rst), .Q(
        \cache[4][2][DATA][23] ) );
  DFFR_X1 \cache_reg[4][2][DATA][22]  ( .D(n286), .CK(net19303), .RN(rst), .Q(
        \cache[4][2][DATA][22] ) );
  DFFR_X1 \cache_reg[4][2][DATA][21]  ( .D(n44), .CK(net19303), .RN(rst), .Q(
        \cache[4][2][DATA][21] ) );
  DFFR_X1 \cache_reg[4][2][DATA][20]  ( .D(n42), .CK(net19303), .RN(rst), .Q(
        \cache[4][2][DATA][20] ) );
  DFFR_X1 \cache_reg[4][2][DATA][19]  ( .D(n48), .CK(net19303), .RN(rst), .Q(
        \cache[4][2][DATA][19] ) );
  DFFR_X1 \cache_reg[4][2][DATA][18]  ( .D(n46), .CK(net19303), .RN(rst), .Q(
        \cache[4][2][DATA][18] ) );
  DFFR_X1 \cache_reg[4][2][DATA][17]  ( .D(n47), .CK(net19303), .RN(rst), .Q(
        \cache[4][2][DATA][17] ) );
  DFFR_X1 \cache_reg[4][2][DATA][16]  ( .D(n279), .CK(net19303), .RN(rst), .Q(
        \cache[4][2][DATA][16] ) );
  DFFR_X1 \cache_reg[4][2][DATA][15]  ( .D(n45), .CK(net19303), .RN(rst), .Q(
        \cache[4][2][DATA][15] ) );
  DFFR_X1 \cache_reg[4][2][DATA][14]  ( .D(n35), .CK(net19303), .RN(n41), .Q(
        \cache[4][2][DATA][14] ) );
  DFFR_X1 \cache_reg[4][2][DATA][13]  ( .D(n52), .CK(net19303), .RN(rst), .Q(
        \cache[4][2][DATA][13] ) );
  DFFR_X1 \cache_reg[4][2][DATA][12]  ( .D(n50), .CK(net19303), .RN(rst), .Q(
        \cache[4][2][DATA][12] ) );
  DFFR_X1 \cache_reg[4][2][DATA][11]  ( .D(n51), .CK(net19303), .RN(rst), .Q(
        \cache[4][2][DATA][11] ) );
  DFFR_X1 \cache_reg[4][2][DATA][10]  ( .D(n49), .CK(net19303), .RN(rst), .Q(
        \cache[4][2][DATA][10] ) );
  DFFR_X1 \cache_reg[4][2][DATA][9]  ( .D(n43), .CK(net19303), .RN(n41), .Q(
        \cache[4][2][DATA][9] ) );
  DFFR_X1 \cache_reg[4][2][DATA][8]  ( .D(n270), .CK(net19303), .RN(n41), .Q(
        \cache[4][2][DATA][8] ) );
  DFFR_X1 \cache_reg[4][2][DATA][7]  ( .D(n204), .CK(net19303), .RN(rst), .Q(
        \cache[4][2][DATA][7] ) );
  DFFR_X1 \cache_reg[4][2][DATA][6]  ( .D(n222), .CK(net19303), .RN(rst), .Q(
        \cache[4][2][DATA][6] ) );
  DFFR_X1 \cache_reg[4][2][DATA][5]  ( .D(n266), .CK(net19303), .RN(rst), .Q(
        \cache[4][2][DATA][5] ) );
  DFFR_X1 \cache_reg[4][2][DATA][4]  ( .D(n264), .CK(net19303), .RN(rst), .Q(
        \cache[4][2][DATA][4] ) );
  DFFR_X1 \cache_reg[4][2][DATA][3]  ( .D(n262), .CK(net19303), .RN(rst), .Q(
        \cache[4][2][DATA][3] ) );
  DFFR_X1 \cache_reg[4][2][DATA][2]  ( .D(n260), .CK(net19303), .RN(rst), .Q(
        \cache[4][2][DATA][2] ) );
  DFFR_X1 \cache_reg[4][2][DATA][1]  ( .D(n216), .CK(net19303), .RN(rst), .Q(
        \cache[4][2][DATA][1] ) );
  DFFR_X1 \cache_reg[4][2][DATA][0]  ( .D(n212), .CK(net19303), .RN(rst), .Q(
        \cache[4][2][DATA][0] ) );
  DFFR_X1 \cache_reg[5][2][DATA][29]  ( .D(n300), .CK(net19363), .RN(rst), .Q(
        \cache[5][2][DATA][29] ) );
  DFFR_X1 \cache_reg[5][2][DATA][28]  ( .D(n298), .CK(net19363), .RN(rst), .Q(
        \cache[5][2][DATA][28] ) );
  DFFR_X1 \cache_reg[5][2][DATA][27]  ( .D(n296), .CK(net19363), .RN(rst), .Q(
        \cache[5][2][DATA][27] ) );
  DFFR_X1 \cache_reg[5][2][DATA][26]  ( .D(n294), .CK(net19363), .RN(rst), .Q(
        \cache[5][2][DATA][26] ) );
  DFFR_X1 \cache_reg[5][2][DATA][25]  ( .D(n292), .CK(net19363), .RN(rst), .Q(
        \cache[5][2][DATA][25] ) );
  DFFR_X1 \cache_reg[5][2][DATA][24]  ( .D(n290), .CK(net19363), .RN(rst), .Q(
        \cache[5][2][DATA][24] ) );
  DFFR_X1 \cache_reg[5][2][DATA][23]  ( .D(n288), .CK(net19363), .RN(rst), .Q(
        \cache[5][2][DATA][23] ) );
  DFFR_X1 \cache_reg[5][2][DATA][22]  ( .D(n286), .CK(net19363), .RN(rst), .Q(
        \cache[5][2][DATA][22] ) );
  DFFR_X1 \cache_reg[5][2][DATA][21]  ( .D(n44), .CK(net19363), .RN(rst), .Q(
        \cache[5][2][DATA][21] ) );
  DFFR_X1 \cache_reg[5][2][DATA][20]  ( .D(n42), .CK(net19363), .RN(rst), .Q(
        \cache[5][2][DATA][20] ) );
  DFFR_X1 \cache_reg[5][2][DATA][19]  ( .D(n48), .CK(net19363), .RN(rst), .Q(
        \cache[5][2][DATA][19] ) );
  DFFR_X1 \cache_reg[5][2][DATA][18]  ( .D(n46), .CK(net19363), .RN(rst), .Q(
        \cache[5][2][DATA][18] ) );
  DFFR_X1 \cache_reg[5][2][DATA][17]  ( .D(n47), .CK(net19363), .RN(rst), .Q(
        \cache[5][2][DATA][17] ) );
  DFFR_X1 \cache_reg[5][2][DATA][16]  ( .D(n279), .CK(net19363), .RN(rst), .Q(
        \cache[5][2][DATA][16] ) );
  DFFR_X1 \cache_reg[5][2][DATA][15]  ( .D(n45), .CK(net19363), .RN(rst), .Q(
        \cache[5][2][DATA][15] ) );
  DFFR_X1 \cache_reg[5][2][DATA][14]  ( .D(n35), .CK(net19363), .RN(rst), .Q(
        \cache[5][2][DATA][14] ) );
  DFFR_X1 \cache_reg[5][2][DATA][13]  ( .D(n52), .CK(net19363), .RN(rst), .Q(
        \cache[5][2][DATA][13] ) );
  DFFR_X1 \cache_reg[5][2][DATA][12]  ( .D(n50), .CK(net19363), .RN(rst), .Q(
        \cache[5][2][DATA][12] ) );
  DFFR_X1 \cache_reg[5][2][DATA][11]  ( .D(n51), .CK(net19363), .RN(n41), .Q(
        \cache[5][2][DATA][11] ) );
  DFFR_X1 \cache_reg[5][2][DATA][10]  ( .D(n49), .CK(net19363), .RN(n41), .Q(
        \cache[5][2][DATA][10] ) );
  DFFR_X1 \cache_reg[5][2][DATA][9]  ( .D(n43), .CK(net19363), .RN(n41), .Q(
        \cache[5][2][DATA][9] ) );
  DFFR_X1 \cache_reg[5][2][DATA][8]  ( .D(n270), .CK(net19363), .RN(n41), .Q(
        \cache[5][2][DATA][8] ) );
  DFFR_X1 \cache_reg[5][2][DATA][7]  ( .D(n204), .CK(net19363), .RN(n41), .Q(
        \cache[5][2][DATA][7] ) );
  DFFR_X1 \cache_reg[5][2][DATA][6]  ( .D(n222), .CK(net19363), .RN(n41), .Q(
        \cache[5][2][DATA][6] ) );
  DFFR_X1 \cache_reg[5][2][DATA][5]  ( .D(n266), .CK(net19363), .RN(n41), .Q(
        \cache[5][2][DATA][5] ) );
  DFFR_X1 \cache_reg[5][2][DATA][4]  ( .D(n264), .CK(net19363), .RN(n41), .Q(
        \cache[5][2][DATA][4] ) );
  DFFR_X1 \cache_reg[5][2][DATA][3]  ( .D(n262), .CK(net19363), .RN(n41), .Q(
        \cache[5][2][DATA][3] ) );
  DFFR_X1 \cache_reg[5][2][DATA][2]  ( .D(n260), .CK(net19363), .RN(n41), .Q(
        \cache[5][2][DATA][2] ) );
  DFFR_X1 \cache_reg[5][2][DATA][1]  ( .D(n216), .CK(net19363), .RN(n41), .Q(
        \cache[5][2][DATA][1] ) );
  DFFR_X1 \cache_reg[5][2][DATA][0]  ( .D(n212), .CK(net19363), .RN(rst), .Q(
        \cache[5][2][DATA][0] ) );
  DFFR_X1 \cache_reg[6][2][DATA][29]  ( .D(n300), .CK(net19423), .RN(n41), .Q(
        \cache[6][2][DATA][29] ) );
  DFFR_X1 \cache_reg[6][2][DATA][28]  ( .D(n298), .CK(net19423), .RN(rst), .Q(
        \cache[6][2][DATA][28] ) );
  DFFR_X1 \cache_reg[6][2][DATA][27]  ( .D(n296), .CK(net19423), .RN(n41), .Q(
        \cache[6][2][DATA][27] ) );
  DFFR_X1 \cache_reg[6][2][DATA][26]  ( .D(n294), .CK(net19423), .RN(n41), .Q(
        \cache[6][2][DATA][26] ) );
  DFFR_X1 \cache_reg[6][2][DATA][25]  ( .D(n292), .CK(net19423), .RN(n41), .Q(
        \cache[6][2][DATA][25] ) );
  DFFR_X1 \cache_reg[6][2][DATA][24]  ( .D(n290), .CK(net19423), .RN(rst), .Q(
        \cache[6][2][DATA][24] ) );
  DFFR_X1 \cache_reg[6][2][DATA][23]  ( .D(n288), .CK(net19423), .RN(rst), .Q(
        \cache[6][2][DATA][23] ) );
  DFFR_X1 \cache_reg[6][2][DATA][22]  ( .D(n286), .CK(net19423), .RN(rst), .Q(
        \cache[6][2][DATA][22] ) );
  DFFR_X1 \cache_reg[6][2][DATA][21]  ( .D(n44), .CK(net19423), .RN(rst), .Q(
        \cache[6][2][DATA][21] ) );
  DFFR_X1 \cache_reg[6][2][DATA][20]  ( .D(n42), .CK(net19423), .RN(n41), .Q(
        \cache[6][2][DATA][20] ) );
  DFFR_X1 \cache_reg[6][2][DATA][19]  ( .D(n48), .CK(net19423), .RN(rst), .Q(
        \cache[6][2][DATA][19] ) );
  DFFR_X1 \cache_reg[6][2][DATA][18]  ( .D(n46), .CK(net19423), .RN(n41), .Q(
        \cache[6][2][DATA][18] ) );
  DFFR_X1 \cache_reg[6][2][DATA][17]  ( .D(n47), .CK(net19423), .RN(rst), .Q(
        \cache[6][2][DATA][17] ) );
  DFFR_X1 \cache_reg[6][2][DATA][16]  ( .D(n279), .CK(net19423), .RN(rst), .Q(
        \cache[6][2][DATA][16] ) );
  DFFR_X1 \cache_reg[6][2][DATA][15]  ( .D(n45), .CK(net19423), .RN(rst), .Q(
        \cache[6][2][DATA][15] ) );
  DFFR_X1 \cache_reg[6][2][DATA][14]  ( .D(n35), .CK(net19423), .RN(rst), .Q(
        \cache[6][2][DATA][14] ) );
  DFFR_X1 \cache_reg[6][2][DATA][13]  ( .D(n52), .CK(net19423), .RN(rst), .Q(
        \cache[6][2][DATA][13] ) );
  DFFR_X1 \cache_reg[6][2][DATA][12]  ( .D(n50), .CK(net19423), .RN(n41), .Q(
        \cache[6][2][DATA][12] ) );
  DFFR_X1 \cache_reg[6][2][DATA][11]  ( .D(n51), .CK(net19423), .RN(rst), .Q(
        \cache[6][2][DATA][11] ) );
  DFFR_X1 \cache_reg[6][2][DATA][10]  ( .D(n49), .CK(net19423), .RN(rst), .Q(
        \cache[6][2][DATA][10] ) );
  DFFR_X1 \cache_reg[6][2][DATA][9]  ( .D(n43), .CK(net19423), .RN(rst), .Q(
        \cache[6][2][DATA][9] ) );
  DFFR_X1 \cache_reg[6][2][DATA][8]  ( .D(n270), .CK(net19423), .RN(rst), .Q(
        \cache[6][2][DATA][8] ) );
  DFFR_X1 \cache_reg[6][2][DATA][7]  ( .D(n204), .CK(net19423), .RN(rst), .Q(
        \cache[6][2][DATA][7] ) );
  DFFR_X1 \cache_reg[6][2][DATA][6]  ( .D(n222), .CK(net19423), .RN(rst), .Q(
        \cache[6][2][DATA][6] ) );
  DFFR_X1 \cache_reg[6][2][DATA][5]  ( .D(n266), .CK(net19423), .RN(rst), .Q(
        \cache[6][2][DATA][5] ) );
  DFFR_X1 \cache_reg[6][2][DATA][4]  ( .D(n264), .CK(net19423), .RN(n41), .Q(
        \cache[6][2][DATA][4] ) );
  DFFR_X1 \cache_reg[6][2][DATA][3]  ( .D(n262), .CK(net19423), .RN(n41), .Q(
        \cache[6][2][DATA][3] ) );
  DFFR_X1 \cache_reg[6][2][DATA][2]  ( .D(n260), .CK(net19423), .RN(n41), .Q(
        \cache[6][2][DATA][2] ) );
  DFFR_X1 \cache_reg[6][2][DATA][1]  ( .D(n216), .CK(net19423), .RN(rst), .Q(
        \cache[6][2][DATA][1] ) );
  DFFR_X1 \cache_reg[6][2][DATA][0]  ( .D(n212), .CK(net19423), .RN(rst), .Q(
        \cache[6][2][DATA][0] ) );
  DFFR_X1 \cache_reg[7][2][DATA][29]  ( .D(n300), .CK(net19483), .RN(n41), .Q(
        \cache[7][2][DATA][29] ) );
  DFFR_X1 \cache_reg[7][2][DATA][28]  ( .D(n298), .CK(net19483), .RN(rst), .Q(
        \cache[7][2][DATA][28] ) );
  DFFR_X1 \cache_reg[7][2][DATA][27]  ( .D(n296), .CK(net19483), .RN(rst), .Q(
        \cache[7][2][DATA][27] ) );
  DFFR_X1 \cache_reg[7][2][DATA][26]  ( .D(n294), .CK(net19483), .RN(rst), .Q(
        \cache[7][2][DATA][26] ) );
  DFFR_X1 \cache_reg[7][2][DATA][25]  ( .D(n292), .CK(net19483), .RN(rst), .Q(
        \cache[7][2][DATA][25] ) );
  DFFR_X1 \cache_reg[7][2][DATA][24]  ( .D(n290), .CK(net19483), .RN(rst), .Q(
        \cache[7][2][DATA][24] ) );
  DFFR_X1 \cache_reg[7][2][DATA][23]  ( .D(n288), .CK(net19483), .RN(n41), .Q(
        \cache[7][2][DATA][23] ) );
  DFFR_X1 \cache_reg[7][2][DATA][22]  ( .D(n286), .CK(net19483), .RN(n41), .Q(
        \cache[7][2][DATA][22] ) );
  DFFR_X1 \cache_reg[7][2][DATA][21]  ( .D(n44), .CK(net19483), .RN(rst), .Q(
        \cache[7][2][DATA][21] ) );
  DFFR_X1 \cache_reg[7][2][DATA][20]  ( .D(n42), .CK(net19483), .RN(rst), .Q(
        \cache[7][2][DATA][20] ) );
  DFFR_X1 \cache_reg[7][2][DATA][19]  ( .D(n48), .CK(net19483), .RN(rst), .Q(
        \cache[7][2][DATA][19] ) );
  DFFR_X1 \cache_reg[7][2][DATA][18]  ( .D(n46), .CK(net19483), .RN(rst), .Q(
        \cache[7][2][DATA][18] ) );
  DFFR_X1 \cache_reg[7][2][DATA][17]  ( .D(n47), .CK(net19483), .RN(rst), .Q(
        \cache[7][2][DATA][17] ) );
  DFFR_X1 \cache_reg[7][2][DATA][16]  ( .D(n279), .CK(net19483), .RN(rst), .Q(
        \cache[7][2][DATA][16] ) );
  DFFR_X1 \cache_reg[7][2][DATA][15]  ( .D(n45), .CK(net19483), .RN(rst), .Q(
        \cache[7][2][DATA][15] ) );
  DFFR_X1 \cache_reg[7][2][DATA][14]  ( .D(n35), .CK(net19483), .RN(rst), .Q(
        \cache[7][2][DATA][14] ) );
  DFFR_X1 \cache_reg[7][2][DATA][13]  ( .D(n52), .CK(net19483), .RN(rst), .Q(
        \cache[7][2][DATA][13] ) );
  DFFR_X1 \cache_reg[7][2][DATA][12]  ( .D(n50), .CK(net19483), .RN(rst), .Q(
        \cache[7][2][DATA][12] ) );
  DFFR_X1 \cache_reg[7][2][DATA][11]  ( .D(n51), .CK(net19483), .RN(rst), .Q(
        \cache[7][2][DATA][11] ) );
  DFFR_X1 \cache_reg[7][2][DATA][10]  ( .D(n49), .CK(net19483), .RN(rst), .Q(
        \cache[7][2][DATA][10] ) );
  DFFR_X1 \cache_reg[7][2][DATA][9]  ( .D(n43), .CK(net19483), .RN(rst), .Q(
        \cache[7][2][DATA][9] ) );
  DFFR_X1 \cache_reg[7][2][DATA][8]  ( .D(n270), .CK(net19483), .RN(rst), .Q(
        \cache[7][2][DATA][8] ) );
  DFFR_X1 \cache_reg[7][2][DATA][7]  ( .D(n204), .CK(net19483), .RN(rst), .Q(
        \cache[7][2][DATA][7] ) );
  DFFR_X1 \cache_reg[7][2][DATA][6]  ( .D(n222), .CK(net19483), .RN(rst), .Q(
        \cache[7][2][DATA][6] ) );
  DFFR_X1 \cache_reg[7][2][DATA][5]  ( .D(n266), .CK(net19483), .RN(rst), .Q(
        \cache[7][2][DATA][5] ) );
  DFFR_X1 \cache_reg[7][2][DATA][4]  ( .D(n264), .CK(net19483), .RN(rst), .Q(
        \cache[7][2][DATA][4] ) );
  DFFR_X1 \cache_reg[7][2][DATA][3]  ( .D(n262), .CK(net19483), .RN(rst), .Q(
        \cache[7][2][DATA][3] ) );
  DFFR_X1 \cache_reg[7][2][DATA][2]  ( .D(n260), .CK(net19483), .RN(rst), .Q(
        \cache[7][2][DATA][2] ) );
  DFFR_X1 \cache_reg[7][2][DATA][1]  ( .D(n216), .CK(net19483), .RN(rst), .Q(
        \cache[7][2][DATA][1] ) );
  DFFR_X1 \cache_reg[7][2][DATA][0]  ( .D(n212), .CK(net19483), .RN(rst), .Q(
        \cache[7][2][DATA][0] ) );
  DFFR_X1 \cache_reg[0][3][DATA][29]  ( .D(n300), .CK(net19078), .RN(rst), .Q(
        \cache[0][3][DATA][29] ) );
  DFFR_X1 \cache_reg[0][3][DATA][28]  ( .D(n298), .CK(net19078), .RN(rst), .Q(
        \cache[0][3][DATA][28] ) );
  DFFR_X1 \cache_reg[0][3][DATA][27]  ( .D(n296), .CK(net19078), .RN(rst), .Q(
        \cache[0][3][DATA][27] ) );
  DFFR_X1 \cache_reg[0][3][DATA][26]  ( .D(n294), .CK(net19078), .RN(rst), .Q(
        \cache[0][3][DATA][26] ) );
  DFFR_X1 \cache_reg[0][3][DATA][25]  ( .D(n292), .CK(net19078), .RN(rst), .Q(
        \cache[0][3][DATA][25] ) );
  DFFR_X1 \cache_reg[0][3][DATA][24]  ( .D(n290), .CK(net19078), .RN(rst), .Q(
        \cache[0][3][DATA][24] ) );
  DFFR_X1 \cache_reg[0][3][DATA][23]  ( .D(n288), .CK(net19078), .RN(rst), .Q(
        \cache[0][3][DATA][23] ) );
  DFFR_X1 \cache_reg[0][3][DATA][22]  ( .D(n286), .CK(net19078), .RN(rst), .Q(
        \cache[0][3][DATA][22] ) );
  DFFR_X1 \cache_reg[0][3][DATA][21]  ( .D(n44), .CK(net19078), .RN(rst), .Q(
        \cache[0][3][DATA][21] ) );
  DFFR_X1 \cache_reg[0][3][DATA][20]  ( .D(n42), .CK(net19078), .RN(rst), .Q(
        \cache[0][3][DATA][20] ) );
  DFFR_X1 \cache_reg[0][3][DATA][19]  ( .D(n48), .CK(net19078), .RN(rst), .Q(
        \cache[0][3][DATA][19] ) );
  DFFR_X1 \cache_reg[0][3][DATA][18]  ( .D(n46), .CK(net19078), .RN(rst), .Q(
        \cache[0][3][DATA][18] ) );
  DFFR_X1 \cache_reg[0][3][DATA][17]  ( .D(n47), .CK(net19078), .RN(rst), .Q(
        \cache[0][3][DATA][17] ) );
  DFFR_X1 \cache_reg[0][3][DATA][16]  ( .D(n279), .CK(net19078), .RN(rst), .Q(
        \cache[0][3][DATA][16] ) );
  DFFR_X1 \cache_reg[0][3][DATA][15]  ( .D(n45), .CK(net19078), .RN(rst), .Q(
        \cache[0][3][DATA][15] ) );
  DFFR_X1 \cache_reg[0][3][DATA][14]  ( .D(n35), .CK(net19078), .RN(rst), .Q(
        \cache[0][3][DATA][14] ) );
  DFFR_X1 \cache_reg[0][3][DATA][13]  ( .D(n52), .CK(net19078), .RN(rst), .Q(
        \cache[0][3][DATA][13] ) );
  DFFR_X1 \cache_reg[0][3][DATA][12]  ( .D(n50), .CK(net19078), .RN(rst), .Q(
        \cache[0][3][DATA][12] ) );
  DFFR_X1 \cache_reg[0][3][DATA][11]  ( .D(n51), .CK(net19078), .RN(rst), .Q(
        \cache[0][3][DATA][11] ) );
  DFFR_X1 \cache_reg[0][3][DATA][10]  ( .D(n49), .CK(net19078), .RN(rst), .Q(
        \cache[0][3][DATA][10] ) );
  DFFR_X1 \cache_reg[0][3][DATA][9]  ( .D(n43), .CK(net19078), .RN(rst), .Q(
        \cache[0][3][DATA][9] ) );
  DFFR_X1 \cache_reg[0][3][DATA][8]  ( .D(n270), .CK(net19078), .RN(rst), .Q(
        \cache[0][3][DATA][8] ) );
  DFFR_X1 \cache_reg[0][3][DATA][7]  ( .D(n204), .CK(net19078), .RN(rst), .Q(
        \cache[0][3][DATA][7] ) );
  DFFR_X1 \cache_reg[0][3][DATA][6]  ( .D(n222), .CK(net19078), .RN(rst), .Q(
        \cache[0][3][DATA][6] ) );
  DFFR_X1 \cache_reg[0][3][DATA][5]  ( .D(n266), .CK(net19078), .RN(rst), .Q(
        \cache[0][3][DATA][5] ) );
  DFFR_X1 \cache_reg[0][3][DATA][4]  ( .D(n264), .CK(net19078), .RN(rst), .Q(
        \cache[0][3][DATA][4] ) );
  DFFR_X1 \cache_reg[0][3][DATA][3]  ( .D(n262), .CK(net19078), .RN(rst), .Q(
        \cache[0][3][DATA][3] ) );
  DFFR_X1 \cache_reg[0][3][DATA][2]  ( .D(n260), .CK(net19078), .RN(rst), .Q(
        \cache[0][3][DATA][2] ) );
  DFFR_X1 \cache_reg[0][3][DATA][1]  ( .D(n216), .CK(net19078), .RN(rst), .Q(
        \cache[0][3][DATA][1] ) );
  DFFR_X1 \cache_reg[0][3][DATA][0]  ( .D(n212), .CK(net19078), .RN(rst), .Q(
        \cache[0][3][DATA][0] ) );
  DFFR_X1 \cache_reg[1][3][DATA][29]  ( .D(n300), .CK(net19138), .RN(rst), .Q(
        \cache[1][3][DATA][29] ) );
  DFFR_X1 \cache_reg[1][3][DATA][28]  ( .D(n298), .CK(net19138), .RN(rst), .Q(
        \cache[1][3][DATA][28] ) );
  DFFR_X1 \cache_reg[1][3][DATA][27]  ( .D(n296), .CK(net19138), .RN(rst), .Q(
        \cache[1][3][DATA][27] ) );
  DFFR_X1 \cache_reg[1][3][DATA][26]  ( .D(n294), .CK(net19138), .RN(rst), .Q(
        \cache[1][3][DATA][26] ) );
  DFFR_X1 \cache_reg[1][3][DATA][25]  ( .D(n292), .CK(net19138), .RN(rst), .Q(
        \cache[1][3][DATA][25] ) );
  DFFR_X1 \cache_reg[1][3][DATA][24]  ( .D(n290), .CK(net19138), .RN(rst), .Q(
        \cache[1][3][DATA][24] ) );
  DFFR_X1 \cache_reg[1][3][DATA][23]  ( .D(n288), .CK(net19138), .RN(rst), .Q(
        \cache[1][3][DATA][23] ) );
  DFFR_X1 \cache_reg[1][3][DATA][22]  ( .D(n286), .CK(net19138), .RN(rst), .Q(
        \cache[1][3][DATA][22] ) );
  DFFR_X1 \cache_reg[1][3][DATA][21]  ( .D(n44), .CK(net19138), .RN(rst), .Q(
        \cache[1][3][DATA][21] ) );
  DFFR_X1 \cache_reg[1][3][DATA][20]  ( .D(n42), .CK(net19138), .RN(rst), .Q(
        \cache[1][3][DATA][20] ) );
  DFFR_X1 \cache_reg[1][3][DATA][19]  ( .D(n48), .CK(net19138), .RN(rst), .Q(
        \cache[1][3][DATA][19] ) );
  DFFR_X1 \cache_reg[1][3][DATA][18]  ( .D(n46), .CK(net19138), .RN(rst), .Q(
        \cache[1][3][DATA][18] ) );
  DFFR_X1 \cache_reg[1][3][DATA][17]  ( .D(n47), .CK(net19138), .RN(rst), .Q(
        \cache[1][3][DATA][17] ) );
  DFFR_X1 \cache_reg[1][3][DATA][16]  ( .D(n279), .CK(net19138), .RN(rst), .Q(
        \cache[1][3][DATA][16] ) );
  DFFR_X1 \cache_reg[1][3][DATA][15]  ( .D(n45), .CK(net19138), .RN(rst), .Q(
        \cache[1][3][DATA][15] ) );
  DFFR_X1 \cache_reg[1][3][DATA][14]  ( .D(n35), .CK(net19138), .RN(rst), .Q(
        \cache[1][3][DATA][14] ) );
  DFFR_X1 \cache_reg[1][3][DATA][13]  ( .D(n52), .CK(net19138), .RN(rst), .Q(
        \cache[1][3][DATA][13] ) );
  DFFR_X1 \cache_reg[1][3][DATA][12]  ( .D(n50), .CK(net19138), .RN(rst), .Q(
        \cache[1][3][DATA][12] ) );
  DFFR_X1 \cache_reg[1][3][DATA][11]  ( .D(n51), .CK(net19138), .RN(rst), .Q(
        \cache[1][3][DATA][11] ) );
  DFFR_X1 \cache_reg[1][3][DATA][10]  ( .D(n49), .CK(net19138), .RN(rst), .Q(
        \cache[1][3][DATA][10] ) );
  DFFR_X1 \cache_reg[1][3][DATA][9]  ( .D(n43), .CK(net19138), .RN(rst), .Q(
        \cache[1][3][DATA][9] ) );
  DFFR_X1 \cache_reg[1][3][DATA][8]  ( .D(n270), .CK(net19138), .RN(rst), .Q(
        \cache[1][3][DATA][8] ) );
  DFFR_X1 \cache_reg[1][3][DATA][7]  ( .D(n204), .CK(net19138), .RN(rst), .Q(
        \cache[1][3][DATA][7] ) );
  DFFR_X1 \cache_reg[1][3][DATA][6]  ( .D(n222), .CK(net19138), .RN(rst), .Q(
        \cache[1][3][DATA][6] ) );
  DFFR_X1 \cache_reg[1][3][DATA][5]  ( .D(n266), .CK(net19138), .RN(rst), .Q(
        \cache[1][3][DATA][5] ) );
  DFFR_X1 \cache_reg[1][3][DATA][4]  ( .D(n264), .CK(net19138), .RN(rst), .Q(
        \cache[1][3][DATA][4] ) );
  DFFR_X1 \cache_reg[1][3][DATA][3]  ( .D(n262), .CK(net19138), .RN(rst), .Q(
        \cache[1][3][DATA][3] ) );
  DFFR_X1 \cache_reg[1][3][DATA][2]  ( .D(n260), .CK(net19138), .RN(rst), .Q(
        \cache[1][3][DATA][2] ) );
  DFFR_X1 \cache_reg[1][3][DATA][1]  ( .D(n216), .CK(net19138), .RN(rst), .Q(
        \cache[1][3][DATA][1] ) );
  DFFR_X1 \cache_reg[1][3][DATA][0]  ( .D(n212), .CK(net19138), .RN(rst), .Q(
        \cache[1][3][DATA][0] ) );
  DFFR_X1 \cache_reg[2][3][DATA][29]  ( .D(n300), .CK(net19198), .RN(rst), .Q(
        \cache[2][3][DATA][29] ) );
  DFFR_X1 \cache_reg[2][3][DATA][28]  ( .D(n298), .CK(net19198), .RN(rst), .Q(
        \cache[2][3][DATA][28] ) );
  DFFR_X1 \cache_reg[2][3][DATA][27]  ( .D(n296), .CK(net19198), .RN(rst), .Q(
        \cache[2][3][DATA][27] ) );
  DFFR_X1 \cache_reg[2][3][DATA][26]  ( .D(n294), .CK(net19198), .RN(rst), .Q(
        \cache[2][3][DATA][26] ) );
  DFFR_X1 \cache_reg[2][3][DATA][25]  ( .D(n292), .CK(net19198), .RN(rst), .Q(
        \cache[2][3][DATA][25] ) );
  DFFR_X1 \cache_reg[2][3][DATA][24]  ( .D(n290), .CK(net19198), .RN(rst), .Q(
        \cache[2][3][DATA][24] ) );
  DFFR_X1 \cache_reg[2][3][DATA][23]  ( .D(n288), .CK(net19198), .RN(rst), .Q(
        \cache[2][3][DATA][23] ) );
  DFFR_X1 \cache_reg[2][3][DATA][22]  ( .D(n286), .CK(net19198), .RN(rst), .Q(
        \cache[2][3][DATA][22] ) );
  DFFR_X1 \cache_reg[2][3][DATA][21]  ( .D(n44), .CK(net19198), .RN(rst), .Q(
        \cache[2][3][DATA][21] ) );
  DFFR_X1 \cache_reg[2][3][DATA][20]  ( .D(n42), .CK(net19198), .RN(rst), .Q(
        \cache[2][3][DATA][20] ) );
  DFFR_X1 \cache_reg[2][3][DATA][19]  ( .D(n48), .CK(net19198), .RN(rst), .Q(
        \cache[2][3][DATA][19] ) );
  DFFR_X1 \cache_reg[2][3][DATA][18]  ( .D(n46), .CK(net19198), .RN(rst), .Q(
        \cache[2][3][DATA][18] ) );
  DFFR_X1 \cache_reg[2][3][DATA][17]  ( .D(n47), .CK(net19198), .RN(rst), .Q(
        \cache[2][3][DATA][17] ) );
  DFFR_X1 \cache_reg[2][3][DATA][16]  ( .D(n279), .CK(net19198), .RN(rst), .Q(
        \cache[2][3][DATA][16] ) );
  DFFR_X1 \cache_reg[2][3][DATA][15]  ( .D(n45), .CK(net19198), .RN(rst), .Q(
        \cache[2][3][DATA][15] ) );
  DFFR_X1 \cache_reg[2][3][DATA][14]  ( .D(n35), .CK(net19198), .RN(rst), .Q(
        \cache[2][3][DATA][14] ) );
  DFFR_X1 \cache_reg[2][3][DATA][13]  ( .D(n52), .CK(net19198), .RN(rst), .Q(
        \cache[2][3][DATA][13] ) );
  DFFR_X1 \cache_reg[2][3][DATA][12]  ( .D(n50), .CK(net19198), .RN(rst), .Q(
        \cache[2][3][DATA][12] ) );
  DFFR_X1 \cache_reg[2][3][DATA][11]  ( .D(n51), .CK(net19198), .RN(rst), .Q(
        \cache[2][3][DATA][11] ) );
  DFFR_X1 \cache_reg[2][3][DATA][10]  ( .D(n49), .CK(net19198), .RN(rst), .Q(
        \cache[2][3][DATA][10] ) );
  DFFR_X1 \cache_reg[2][3][DATA][9]  ( .D(n43), .CK(net19198), .RN(rst), .Q(
        \cache[2][3][DATA][9] ) );
  DFFR_X1 \cache_reg[2][3][DATA][8]  ( .D(n270), .CK(net19198), .RN(rst), .Q(
        \cache[2][3][DATA][8] ) );
  DFFR_X1 \cache_reg[2][3][DATA][7]  ( .D(n204), .CK(net19198), .RN(rst), .Q(
        \cache[2][3][DATA][7] ) );
  DFFR_X1 \cache_reg[2][3][DATA][6]  ( .D(n222), .CK(net19198), .RN(rst), .Q(
        \cache[2][3][DATA][6] ) );
  DFFR_X1 \cache_reg[2][3][DATA][5]  ( .D(n266), .CK(net19198), .RN(rst), .Q(
        \cache[2][3][DATA][5] ) );
  DFFR_X1 \cache_reg[2][3][DATA][4]  ( .D(n264), .CK(net19198), .RN(rst), .Q(
        \cache[2][3][DATA][4] ) );
  DFFR_X1 \cache_reg[2][3][DATA][3]  ( .D(n262), .CK(net19198), .RN(rst), .Q(
        \cache[2][3][DATA][3] ) );
  DFFR_X1 \cache_reg[2][3][DATA][2]  ( .D(n260), .CK(net19198), .RN(rst), .Q(
        \cache[2][3][DATA][2] ) );
  DFFR_X1 \cache_reg[2][3][DATA][1]  ( .D(n216), .CK(net19198), .RN(rst), .Q(
        \cache[2][3][DATA][1] ) );
  DFFR_X1 \cache_reg[2][3][DATA][0]  ( .D(n212), .CK(net19198), .RN(rst), .Q(
        \cache[2][3][DATA][0] ) );
  DFFR_X1 \cache_reg[3][3][DATA][29]  ( .D(n300), .CK(net19258), .RN(rst), .Q(
        \cache[3][3][DATA][29] ) );
  DFFR_X1 \cache_reg[3][3][DATA][28]  ( .D(n298), .CK(net19258), .RN(rst), .Q(
        \cache[3][3][DATA][28] ) );
  DFFR_X1 \cache_reg[3][3][DATA][27]  ( .D(n296), .CK(net19258), .RN(rst), .Q(
        \cache[3][3][DATA][27] ) );
  DFFR_X1 \cache_reg[3][3][DATA][26]  ( .D(n294), .CK(net19258), .RN(rst), .Q(
        \cache[3][3][DATA][26] ) );
  DFFR_X1 \cache_reg[3][3][DATA][25]  ( .D(n292), .CK(net19258), .RN(rst), .Q(
        \cache[3][3][DATA][25] ) );
  DFFR_X1 \cache_reg[3][3][DATA][24]  ( .D(n290), .CK(net19258), .RN(rst), .Q(
        \cache[3][3][DATA][24] ) );
  DFFR_X1 \cache_reg[3][3][DATA][23]  ( .D(n288), .CK(net19258), .RN(n304), 
        .Q(\cache[3][3][DATA][23] ) );
  DFFR_X1 \cache_reg[3][3][DATA][22]  ( .D(n286), .CK(net19258), .RN(rst), .Q(
        \cache[3][3][DATA][22] ) );
  DFFR_X1 \cache_reg[3][3][DATA][21]  ( .D(n44), .CK(net19258), .RN(rst), .Q(
        \cache[3][3][DATA][21] ) );
  DFFR_X1 \cache_reg[3][3][DATA][20]  ( .D(n42), .CK(net19258), .RN(rst), .Q(
        \cache[3][3][DATA][20] ) );
  DFFR_X1 \cache_reg[3][3][DATA][19]  ( .D(n48), .CK(net19258), .RN(rst), .Q(
        \cache[3][3][DATA][19] ) );
  DFFR_X1 \cache_reg[3][3][DATA][18]  ( .D(n46), .CK(net19258), .RN(rst), .Q(
        \cache[3][3][DATA][18] ) );
  DFFR_X1 \cache_reg[3][3][DATA][17]  ( .D(n47), .CK(net19258), .RN(rst), .Q(
        \cache[3][3][DATA][17] ) );
  DFFR_X1 \cache_reg[3][3][DATA][16]  ( .D(n279), .CK(net19258), .RN(rst), .Q(
        \cache[3][3][DATA][16] ) );
  DFFR_X1 \cache_reg[3][3][DATA][15]  ( .D(n45), .CK(net19258), .RN(rst), .Q(
        \cache[3][3][DATA][15] ) );
  DFFR_X1 \cache_reg[3][3][DATA][14]  ( .D(n35), .CK(net19258), .RN(rst), .Q(
        \cache[3][3][DATA][14] ) );
  DFFR_X1 \cache_reg[3][3][DATA][13]  ( .D(n52), .CK(net19258), .RN(rst), .Q(
        \cache[3][3][DATA][13] ) );
  DFFR_X1 \cache_reg[3][3][DATA][12]  ( .D(n50), .CK(net19258), .RN(rst), .Q(
        \cache[3][3][DATA][12] ) );
  DFFR_X1 \cache_reg[3][3][DATA][11]  ( .D(n51), .CK(net19258), .RN(rst), .Q(
        \cache[3][3][DATA][11] ) );
  DFFR_X1 \cache_reg[3][3][DATA][10]  ( .D(n49), .CK(net19258), .RN(rst), .Q(
        \cache[3][3][DATA][10] ) );
  DFFR_X1 \cache_reg[3][3][DATA][9]  ( .D(n43), .CK(net19258), .RN(n304), .Q(
        \cache[3][3][DATA][9] ) );
  DFFR_X1 \cache_reg[3][3][DATA][8]  ( .D(n270), .CK(net19258), .RN(rst), .Q(
        \cache[3][3][DATA][8] ) );
  DFFR_X1 \cache_reg[3][3][DATA][7]  ( .D(n204), .CK(net19258), .RN(rst), .Q(
        \cache[3][3][DATA][7] ) );
  DFFR_X1 \cache_reg[3][3][DATA][6]  ( .D(n222), .CK(net19258), .RN(rst), .Q(
        \cache[3][3][DATA][6] ) );
  DFFR_X1 \cache_reg[3][3][DATA][5]  ( .D(n266), .CK(net19258), .RN(rst), .Q(
        \cache[3][3][DATA][5] ) );
  DFFR_X1 \cache_reg[3][3][DATA][4]  ( .D(n264), .CK(net19258), .RN(rst), .Q(
        \cache[3][3][DATA][4] ) );
  DFFR_X1 \cache_reg[3][3][DATA][3]  ( .D(n262), .CK(net19258), .RN(rst), .Q(
        \cache[3][3][DATA][3] ) );
  DFFR_X1 \cache_reg[3][3][DATA][2]  ( .D(n260), .CK(net19258), .RN(rst), .Q(
        \cache[3][3][DATA][2] ) );
  DFFR_X1 \cache_reg[3][3][DATA][1]  ( .D(n216), .CK(net19258), .RN(rst), .Q(
        \cache[3][3][DATA][1] ) );
  DFFR_X1 \cache_reg[3][3][DATA][0]  ( .D(n212), .CK(net19258), .RN(rst), .Q(
        \cache[3][3][DATA][0] ) );
  DFFR_X1 \cache_reg[4][3][DATA][29]  ( .D(n300), .CK(net19318), .RN(rst), .Q(
        \cache[4][3][DATA][29] ) );
  DFFR_X1 \cache_reg[4][3][DATA][28]  ( .D(n298), .CK(net19318), .RN(n304), 
        .Q(\cache[4][3][DATA][28] ) );
  DFFR_X1 \cache_reg[4][3][DATA][27]  ( .D(n296), .CK(net19318), .RN(rst), .Q(
        \cache[4][3][DATA][27] ) );
  DFFR_X1 \cache_reg[4][3][DATA][26]  ( .D(n294), .CK(net19318), .RN(rst), .Q(
        \cache[4][3][DATA][26] ) );
  DFFR_X1 \cache_reg[4][3][DATA][25]  ( .D(n292), .CK(net19318), .RN(rst), .Q(
        \cache[4][3][DATA][25] ) );
  DFFR_X1 \cache_reg[4][3][DATA][24]  ( .D(n290), .CK(net19318), .RN(rst), .Q(
        \cache[4][3][DATA][24] ) );
  DFFR_X1 \cache_reg[4][3][DATA][23]  ( .D(n288), .CK(net19318), .RN(rst), .Q(
        \cache[4][3][DATA][23] ) );
  DFFR_X1 \cache_reg[4][3][DATA][22]  ( .D(n286), .CK(net19318), .RN(rst), .Q(
        \cache[4][3][DATA][22] ) );
  DFFR_X1 \cache_reg[4][3][DATA][21]  ( .D(n44), .CK(net19318), .RN(rst), .Q(
        \cache[4][3][DATA][21] ) );
  DFFR_X1 \cache_reg[4][3][DATA][20]  ( .D(n42), .CK(net19318), .RN(rst), .Q(
        \cache[4][3][DATA][20] ) );
  DFFR_X1 \cache_reg[4][3][DATA][19]  ( .D(n48), .CK(net19318), .RN(rst), .Q(
        \cache[4][3][DATA][19] ) );
  DFFR_X1 \cache_reg[4][3][DATA][18]  ( .D(n46), .CK(net19318), .RN(rst), .Q(
        \cache[4][3][DATA][18] ) );
  DFFR_X1 \cache_reg[4][3][DATA][17]  ( .D(n47), .CK(net19318), .RN(rst), .Q(
        \cache[4][3][DATA][17] ) );
  DFFR_X1 \cache_reg[4][3][DATA][16]  ( .D(n279), .CK(net19318), .RN(rst), .Q(
        \cache[4][3][DATA][16] ) );
  DFFR_X1 \cache_reg[4][3][DATA][15]  ( .D(n45), .CK(net19318), .RN(rst), .Q(
        \cache[4][3][DATA][15] ) );
  DFFR_X1 \cache_reg[4][3][DATA][14]  ( .D(n35), .CK(net19318), .RN(rst), .Q(
        \cache[4][3][DATA][14] ) );
  DFFR_X1 \cache_reg[4][3][DATA][13]  ( .D(n52), .CK(net19318), .RN(rst), .Q(
        \cache[4][3][DATA][13] ) );
  DFFR_X1 \cache_reg[4][3][DATA][12]  ( .D(n50), .CK(net19318), .RN(rst), .Q(
        \cache[4][3][DATA][12] ) );
  DFFR_X1 \cache_reg[4][3][DATA][11]  ( .D(n51), .CK(net19318), .RN(rst), .Q(
        \cache[4][3][DATA][11] ) );
  DFFR_X1 \cache_reg[4][3][DATA][10]  ( .D(n49), .CK(net19318), .RN(rst), .Q(
        \cache[4][3][DATA][10] ) );
  DFFR_X1 \cache_reg[4][3][DATA][9]  ( .D(n43), .CK(net19318), .RN(rst), .Q(
        \cache[4][3][DATA][9] ) );
  DFFR_X1 \cache_reg[4][3][DATA][8]  ( .D(n270), .CK(net19318), .RN(rst), .Q(
        \cache[4][3][DATA][8] ) );
  DFFR_X1 \cache_reg[4][3][DATA][7]  ( .D(n204), .CK(net19318), .RN(rst), .Q(
        \cache[4][3][DATA][7] ) );
  DFFR_X1 \cache_reg[4][3][DATA][6]  ( .D(n222), .CK(net19318), .RN(rst), .Q(
        \cache[4][3][DATA][6] ) );
  DFFR_X1 \cache_reg[4][3][DATA][5]  ( .D(n266), .CK(net19318), .RN(rst), .Q(
        \cache[4][3][DATA][5] ) );
  DFFR_X1 \cache_reg[4][3][DATA][4]  ( .D(n264), .CK(net19318), .RN(rst), .Q(
        \cache[4][3][DATA][4] ) );
  DFFR_X1 \cache_reg[4][3][DATA][3]  ( .D(n262), .CK(net19318), .RN(rst), .Q(
        \cache[4][3][DATA][3] ) );
  DFFR_X1 \cache_reg[4][3][DATA][2]  ( .D(n260), .CK(net19318), .RN(rst), .Q(
        \cache[4][3][DATA][2] ) );
  DFFR_X1 \cache_reg[4][3][DATA][1]  ( .D(n216), .CK(net19318), .RN(rst), .Q(
        \cache[4][3][DATA][1] ) );
  DFFR_X1 \cache_reg[4][3][DATA][0]  ( .D(n212), .CK(net19318), .RN(rst), .Q(
        \cache[4][3][DATA][0] ) );
  DFFR_X1 \cache_reg[5][3][DATA][29]  ( .D(n300), .CK(net19378), .RN(rst), .Q(
        \cache[5][3][DATA][29] ) );
  DFFR_X1 \cache_reg[5][3][DATA][28]  ( .D(n298), .CK(net19378), .RN(rst), .Q(
        \cache[5][3][DATA][28] ) );
  DFFR_X1 \cache_reg[5][3][DATA][27]  ( .D(n296), .CK(net19378), .RN(rst), .Q(
        \cache[5][3][DATA][27] ) );
  DFFR_X1 \cache_reg[5][3][DATA][26]  ( .D(n294), .CK(net19378), .RN(rst), .Q(
        \cache[5][3][DATA][26] ) );
  DFFR_X1 \cache_reg[5][3][DATA][25]  ( .D(n292), .CK(net19378), .RN(rst), .Q(
        \cache[5][3][DATA][25] ) );
  DFFR_X1 \cache_reg[5][3][DATA][24]  ( .D(n290), .CK(net19378), .RN(rst), .Q(
        \cache[5][3][DATA][24] ) );
  DFFR_X1 \cache_reg[5][3][DATA][23]  ( .D(n288), .CK(net19378), .RN(rst), .Q(
        \cache[5][3][DATA][23] ) );
  DFFR_X1 \cache_reg[5][3][DATA][22]  ( .D(n286), .CK(net19378), .RN(rst), .Q(
        \cache[5][3][DATA][22] ) );
  DFFR_X1 \cache_reg[5][3][DATA][21]  ( .D(n44), .CK(net19378), .RN(rst), .Q(
        \cache[5][3][DATA][21] ) );
  DFFR_X1 \cache_reg[5][3][DATA][20]  ( .D(n42), .CK(net19378), .RN(rst), .Q(
        \cache[5][3][DATA][20] ) );
  DFFR_X1 \cache_reg[5][3][DATA][19]  ( .D(n48), .CK(net19378), .RN(rst), .Q(
        \cache[5][3][DATA][19] ) );
  DFFR_X1 \cache_reg[5][3][DATA][18]  ( .D(n46), .CK(net19378), .RN(rst), .Q(
        \cache[5][3][DATA][18] ) );
  DFFR_X1 \cache_reg[5][3][DATA][17]  ( .D(n47), .CK(net19378), .RN(rst), .Q(
        \cache[5][3][DATA][17] ) );
  DFFR_X1 \cache_reg[5][3][DATA][16]  ( .D(n279), .CK(net19378), .RN(rst), .Q(
        \cache[5][3][DATA][16] ) );
  DFFR_X1 \cache_reg[5][3][DATA][15]  ( .D(n45), .CK(net19378), .RN(rst), .Q(
        \cache[5][3][DATA][15] ) );
  DFFR_X1 \cache_reg[5][3][DATA][14]  ( .D(n35), .CK(net19378), .RN(rst), .Q(
        \cache[5][3][DATA][14] ) );
  DFFR_X1 \cache_reg[5][3][DATA][13]  ( .D(n52), .CK(net19378), .RN(rst), .Q(
        \cache[5][3][DATA][13] ) );
  DFFR_X1 \cache_reg[5][3][DATA][12]  ( .D(n50), .CK(net19378), .RN(rst), .Q(
        \cache[5][3][DATA][12] ) );
  DFFR_X1 \cache_reg[5][3][DATA][11]  ( .D(n51), .CK(net19378), .RN(rst), .Q(
        \cache[5][3][DATA][11] ) );
  DFFR_X1 \cache_reg[5][3][DATA][10]  ( .D(n49), .CK(net19378), .RN(rst), .Q(
        \cache[5][3][DATA][10] ) );
  DFFR_X1 \cache_reg[5][3][DATA][9]  ( .D(n43), .CK(net19378), .RN(rst), .Q(
        \cache[5][3][DATA][9] ) );
  DFFR_X1 \cache_reg[5][3][DATA][8]  ( .D(n270), .CK(net19378), .RN(rst), .Q(
        \cache[5][3][DATA][8] ) );
  DFFR_X1 \cache_reg[5][3][DATA][7]  ( .D(n204), .CK(net19378), .RN(rst), .Q(
        \cache[5][3][DATA][7] ) );
  DFFR_X1 \cache_reg[5][3][DATA][6]  ( .D(n222), .CK(net19378), .RN(rst), .Q(
        \cache[5][3][DATA][6] ) );
  DFFR_X1 \cache_reg[5][3][DATA][5]  ( .D(n266), .CK(net19378), .RN(rst), .Q(
        \cache[5][3][DATA][5] ) );
  DFFR_X1 \cache_reg[5][3][DATA][4]  ( .D(n264), .CK(net19378), .RN(rst), .Q(
        \cache[5][3][DATA][4] ) );
  DFFR_X1 \cache_reg[5][3][DATA][3]  ( .D(n262), .CK(net19378), .RN(rst), .Q(
        \cache[5][3][DATA][3] ) );
  DFFR_X1 \cache_reg[5][3][DATA][2]  ( .D(n260), .CK(net19378), .RN(n304), .Q(
        \cache[5][3][DATA][2] ) );
  DFFR_X1 \cache_reg[5][3][DATA][1]  ( .D(n216), .CK(net19378), .RN(rst), .Q(
        \cache[5][3][DATA][1] ) );
  DFFR_X1 \cache_reg[5][3][DATA][0]  ( .D(n212), .CK(net19378), .RN(n304), .Q(
        \cache[5][3][DATA][0] ) );
  DFFR_X1 \cache_reg[6][3][DATA][29]  ( .D(n300), .CK(net19438), .RN(rst), .Q(
        \cache[6][3][DATA][29] ) );
  DFFR_X1 \cache_reg[6][3][DATA][28]  ( .D(n298), .CK(net19438), .RN(rst), .Q(
        \cache[6][3][DATA][28] ) );
  DFFR_X1 \cache_reg[6][3][DATA][27]  ( .D(n296), .CK(net19438), .RN(rst), .Q(
        \cache[6][3][DATA][27] ) );
  DFFR_X1 \cache_reg[6][3][DATA][26]  ( .D(n294), .CK(net19438), .RN(rst), .Q(
        \cache[6][3][DATA][26] ) );
  DFFR_X1 \cache_reg[6][3][DATA][25]  ( .D(n292), .CK(net19438), .RN(rst), .Q(
        \cache[6][3][DATA][25] ) );
  DFFR_X1 \cache_reg[6][3][DATA][24]  ( .D(n290), .CK(net19438), .RN(rst), .Q(
        \cache[6][3][DATA][24] ) );
  DFFR_X1 \cache_reg[6][3][DATA][23]  ( .D(n288), .CK(net19438), .RN(rst), .Q(
        \cache[6][3][DATA][23] ) );
  DFFR_X1 \cache_reg[6][3][DATA][22]  ( .D(n286), .CK(net19438), .RN(n304), 
        .Q(\cache[6][3][DATA][22] ) );
  DFFR_X1 \cache_reg[6][3][DATA][21]  ( .D(n44), .CK(net19438), .RN(rst), .Q(
        \cache[6][3][DATA][21] ) );
  DFFR_X1 \cache_reg[6][3][DATA][20]  ( .D(n42), .CK(net19438), .RN(rst), .Q(
        \cache[6][3][DATA][20] ) );
  DFFR_X1 \cache_reg[6][3][DATA][19]  ( .D(n48), .CK(net19438), .RN(rst), .Q(
        \cache[6][3][DATA][19] ) );
  DFFR_X1 \cache_reg[6][3][DATA][18]  ( .D(n46), .CK(net19438), .RN(rst), .Q(
        \cache[6][3][DATA][18] ) );
  DFFR_X1 \cache_reg[6][3][DATA][17]  ( .D(n47), .CK(net19438), .RN(rst), .Q(
        \cache[6][3][DATA][17] ) );
  DFFR_X1 \cache_reg[6][3][DATA][16]  ( .D(n279), .CK(net19438), .RN(rst), .Q(
        \cache[6][3][DATA][16] ) );
  DFFR_X1 \cache_reg[6][3][DATA][15]  ( .D(n45), .CK(net19438), .RN(n304), .Q(
        \cache[6][3][DATA][15] ) );
  DFFR_X1 \cache_reg[6][3][DATA][14]  ( .D(n35), .CK(net19438), .RN(rst), .Q(
        \cache[6][3][DATA][14] ) );
  DFFR_X1 \cache_reg[6][3][DATA][13]  ( .D(n52), .CK(net19438), .RN(rst), .Q(
        \cache[6][3][DATA][13] ) );
  DFFR_X1 \cache_reg[6][3][DATA][12]  ( .D(n50), .CK(net19438), .RN(rst), .Q(
        \cache[6][3][DATA][12] ) );
  DFFR_X1 \cache_reg[6][3][DATA][11]  ( .D(n51), .CK(net19438), .RN(rst), .Q(
        \cache[6][3][DATA][11] ) );
  DFFR_X1 \cache_reg[6][3][DATA][10]  ( .D(n49), .CK(net19438), .RN(rst), .Q(
        \cache[6][3][DATA][10] ) );
  DFFR_X1 \cache_reg[6][3][DATA][9]  ( .D(n43), .CK(net19438), .RN(rst), .Q(
        \cache[6][3][DATA][9] ) );
  DFFR_X1 \cache_reg[6][3][DATA][8]  ( .D(n270), .CK(net19438), .RN(rst), .Q(
        \cache[6][3][DATA][8] ) );
  DFFR_X1 \cache_reg[6][3][DATA][7]  ( .D(n204), .CK(net19438), .RN(rst), .Q(
        \cache[6][3][DATA][7] ) );
  DFFR_X1 \cache_reg[6][3][DATA][6]  ( .D(n222), .CK(net19438), .RN(rst), .Q(
        \cache[6][3][DATA][6] ) );
  DFFR_X1 \cache_reg[6][3][DATA][5]  ( .D(n266), .CK(net19438), .RN(rst), .Q(
        \cache[6][3][DATA][5] ) );
  DFFR_X1 \cache_reg[6][3][DATA][4]  ( .D(n264), .CK(net19438), .RN(rst), .Q(
        \cache[6][3][DATA][4] ) );
  DFFR_X1 \cache_reg[6][3][DATA][3]  ( .D(n262), .CK(net19438), .RN(rst), .Q(
        \cache[6][3][DATA][3] ) );
  DFFR_X1 \cache_reg[6][3][DATA][2]  ( .D(n260), .CK(net19438), .RN(n304), .Q(
        \cache[6][3][DATA][2] ) );
  DFFR_X1 \cache_reg[6][3][DATA][1]  ( .D(n216), .CK(net19438), .RN(rst), .Q(
        \cache[6][3][DATA][1] ) );
  DFFR_X1 \cache_reg[6][3][DATA][0]  ( .D(n212), .CK(net19438), .RN(rst), .Q(
        \cache[6][3][DATA][0] ) );
  DFFR_X1 \cache_reg[7][3][DATA][29]  ( .D(n300), .CK(net19498), .RN(rst), .Q(
        \cache[7][3][DATA][29] ) );
  DFFR_X1 \cache_reg[7][3][DATA][28]  ( .D(n298), .CK(net19498), .RN(rst), .Q(
        \cache[7][3][DATA][28] ) );
  DFFR_X1 \cache_reg[7][3][DATA][27]  ( .D(n296), .CK(net19498), .RN(rst), .Q(
        \cache[7][3][DATA][27] ) );
  DFFR_X1 \cache_reg[7][3][DATA][26]  ( .D(n294), .CK(net19498), .RN(rst), .Q(
        \cache[7][3][DATA][26] ) );
  DFFR_X1 \cache_reg[7][3][DATA][25]  ( .D(n292), .CK(net19498), .RN(n304), 
        .Q(\cache[7][3][DATA][25] ) );
  DFFR_X1 \cache_reg[7][3][DATA][24]  ( .D(n290), .CK(net19498), .RN(rst), .Q(
        \cache[7][3][DATA][24] ) );
  DFFR_X1 \cache_reg[7][3][DATA][23]  ( .D(n288), .CK(net19498), .RN(rst), .Q(
        \cache[7][3][DATA][23] ) );
  DFFR_X1 \cache_reg[7][3][DATA][22]  ( .D(n286), .CK(net19498), .RN(n304), 
        .Q(\cache[7][3][DATA][22] ) );
  DFFR_X1 \cache_reg[7][3][DATA][21]  ( .D(n44), .CK(net19498), .RN(rst), .Q(
        \cache[7][3][DATA][21] ) );
  DFFR_X1 \cache_reg[7][3][DATA][20]  ( .D(n42), .CK(net19498), .RN(rst), .Q(
        \cache[7][3][DATA][20] ) );
  DFFR_X1 \cache_reg[7][3][DATA][19]  ( .D(n48), .CK(net19498), .RN(rst), .Q(
        \cache[7][3][DATA][19] ) );
  DFFR_X1 \cache_reg[7][3][DATA][18]  ( .D(n46), .CK(net19498), .RN(rst), .Q(
        \cache[7][3][DATA][18] ) );
  DFFR_X1 \cache_reg[7][3][DATA][17]  ( .D(n47), .CK(net19498), .RN(rst), .Q(
        \cache[7][3][DATA][17] ) );
  DFFR_X1 \cache_reg[7][3][DATA][16]  ( .D(n279), .CK(net19498), .RN(rst), .Q(
        \cache[7][3][DATA][16] ) );
  DFFR_X1 \cache_reg[7][3][DATA][15]  ( .D(n45), .CK(net19498), .RN(rst), .Q(
        \cache[7][3][DATA][15] ) );
  DFFR_X1 \cache_reg[7][3][DATA][14]  ( .D(n35), .CK(net19498), .RN(rst), .Q(
        \cache[7][3][DATA][14] ) );
  DFFR_X1 \cache_reg[7][3][DATA][13]  ( .D(n52), .CK(net19498), .RN(n304), .Q(
        \cache[7][3][DATA][13] ) );
  DFFR_X1 \cache_reg[7][3][DATA][12]  ( .D(n50), .CK(net19498), .RN(rst), .Q(
        \cache[7][3][DATA][12] ) );
  DFFR_X1 \cache_reg[7][3][DATA][11]  ( .D(n51), .CK(net19498), .RN(rst), .Q(
        \cache[7][3][DATA][11] ) );
  DFFR_X1 \cache_reg[7][3][DATA][10]  ( .D(n49), .CK(net19498), .RN(rst), .Q(
        \cache[7][3][DATA][10] ) );
  DFFR_X1 \cache_reg[7][3][DATA][9]  ( .D(n43), .CK(net19498), .RN(n304), .Q(
        \cache[7][3][DATA][9] ) );
  DFFR_X1 \cache_reg[7][3][DATA][8]  ( .D(n270), .CK(net19498), .RN(n304), .Q(
        \cache[7][3][DATA][8] ) );
  DFFR_X1 \cache_reg[7][3][DATA][7]  ( .D(n204), .CK(net19498), .RN(rst), .Q(
        \cache[7][3][DATA][7] ) );
  DFFR_X1 \cache_reg[7][3][DATA][6]  ( .D(n222), .CK(net19498), .RN(n304), .Q(
        \cache[7][3][DATA][6] ) );
  DFFR_X1 \cache_reg[7][3][DATA][5]  ( .D(n266), .CK(net19498), .RN(rst), .Q(
        \cache[7][3][DATA][5] ) );
  DFFR_X1 \cache_reg[7][3][DATA][4]  ( .D(n264), .CK(net19498), .RN(rst), .Q(
        \cache[7][3][DATA][4] ) );
  DFFR_X1 \cache_reg[7][3][DATA][3]  ( .D(n262), .CK(net19498), .RN(rst), .Q(
        \cache[7][3][DATA][3] ) );
  DFFR_X1 \cache_reg[7][3][DATA][2]  ( .D(n260), .CK(net19498), .RN(rst), .Q(
        \cache[7][3][DATA][2] ) );
  DFFR_X1 \cache_reg[7][3][DATA][1]  ( .D(n216), .CK(net19498), .RN(rst), .Q(
        \cache[7][3][DATA][1] ) );
  DFFR_X1 \cache_reg[7][3][DATA][0]  ( .D(n212), .CK(net19498), .RN(rst), .Q(
        \cache[7][3][DATA][0] ) );
  DFFS_X1 \last_prediction_reg[2]  ( .D(n27), .CK(net19518), .SN(rst), .Q(n110) );
  DFFR_X1 \last_prediction_reg[9]  ( .D(pc_out[9]), .CK(net19513), .RN(rst), 
        .QN(n124) );
  DFFR_X1 \last_prediction_reg[8]  ( .D(pc_out[8]), .CK(net19518), .RN(rst), 
        .QN(n123) );
  DFFR_X1 \last_prediction_reg[3]  ( .D(pc_out[3]), .CK(net19518), .RN(rst), 
        .QN(n111) );
  DFFR_X1 \last_prediction_reg[16]  ( .D(pc_out[16]), .CK(net19513), .RN(n304), 
        .QN(n117) );
  DFFS_X1 \last_set_reg[0]  ( .D(n609), .CK(net19518), .SN(rst), .Q(n119), 
        .QN(\last_set[0] ) );
  DFFS_X1 \last_set_reg[1]  ( .D(pc_fetch[3]), .CK(net19518), .SN(rst), .Q(
        n105), .QN(\last_set[1] ) );
  DFFS_X1 verify_reg ( .D(n606), .CK(net19508), .SN(rst), .Q(n108), .QN(verify) );
  DFFR_X1 \last_prediction_reg[25]  ( .D(pc_out[25]), .CK(net19513), .RN(rst), 
        .Q(last_prediction[25]), .QN(n116) );
  DFFR_X1 \last_prediction_reg[23]  ( .D(pc_out[23]), .CK(net19513), .RN(rst), 
        .Q(last_prediction[23]), .QN(n139) );
  DFFR_X1 \last_prediction_reg[20]  ( .D(pc_out[20]), .CK(net19513), .RN(n304), 
        .QN(n74) );
  DFFR_X1 \last_prediction_reg[19]  ( .D(pc_out[19]), .CK(net19513), .RN(n304), 
        .QN(n75) );
  DFFR_X1 \last_prediction_reg[18]  ( .D(pc_out[18]), .CK(net19513), .RN(n304), 
        .QN(n77) );
  DFFR_X1 \last_prediction_reg[14]  ( .D(pc_out[14]), .CK(net19513), .RN(n304), 
        .Q(last_prediction[14]), .QN(n113) );
  DFFR_X1 \last_prediction_reg[15]  ( .D(pc_out[15]), .CK(net19513), .RN(n304), 
        .Q(last_prediction[15]), .QN(n126) );
  DFFR_X1 \last_prediction_reg[17]  ( .D(pc_out[17]), .CK(net19513), .RN(n304), 
        .QN(n79) );
  DFFR_X1 \last_prediction_reg[11]  ( .D(pc_out[11]), .CK(net19513), .RN(n304), 
        .Q(last_prediction[11]), .QN(n114) );
  DFFR_X1 \last_prediction_reg[13]  ( .D(pc_out[13]), .CK(net19513), .RN(n304), 
        .Q(last_prediction[13]), .QN(n125) );
  DFFR_X1 \last_prediction_reg[12]  ( .D(pc_out[12]), .CK(net19513), .RN(n304), 
        .Q(last_prediction[12]), .QN(n112) );
  DFFR_X1 \last_prediction_reg[10]  ( .D(pc_out[10]), .CK(net19513), .RN(rst), 
        .Q(last_prediction[10]), .QN(n135) );
  DFFR_X1 \last_prediction_reg[24]  ( .D(pc_out[24]), .CK(net19513), .RN(rst), 
        .Q(last_prediction[24]), .QN(n137) );
  DFFR_X1 \last_prediction_reg[7]  ( .D(pc_out[7]), .CK(net19518), .RN(rst), 
        .Q(last_prediction[7]), .QN(n133) );
  DFFR_X1 \last_prediction_reg[5]  ( .D(pc_out[5]), .CK(net19518), .RN(rst), 
        .Q(last_prediction[5]), .QN(n115) );
  DFFR_X1 \last_prediction_reg[27]  ( .D(pc_out[27]), .CK(net19513), .RN(rst), 
        .Q(last_prediction[27]), .QN(n134) );
  DFFR_X1 \last_prediction_reg[22]  ( .D(pc_out[22]), .CK(net19513), .RN(rst), 
        .QN(n73) );
  DFFR_X1 \last_prediction_reg[21]  ( .D(pc_out[21]), .CK(net19513), .RN(n304), 
        .Q(last_prediction[21]), .QN(n138) );
  DFFR_X1 \last_prediction_reg[30]  ( .D(pc_out[30]), .CK(net19513), .RN(rst), 
        .Q(last_prediction[30]), .QN(n128) );
  DFFR_X1 \last_prediction_reg[28]  ( .D(pc_out[28]), .CK(net19513), .RN(rst), 
        .Q(last_prediction[28]), .QN(n127) );
  DFFR_X1 \last_prediction_reg[26]  ( .D(pc_out[26]), .CK(net19513), .RN(rst), 
        .Q(last_prediction[26]), .QN(n130) );
  DFFR_X1 \last_prediction_reg[31]  ( .D(pc_out[31]), .CK(net19513), .RN(rst), 
        .Q(last_prediction[31]), .QN(n132) );
  DFFR_X1 \last_prediction_reg[4]  ( .D(pc_out[4]), .CK(net19518), .RN(rst), 
        .Q(last_prediction[4]), .QN(n136) );
  DFFR_X1 \last_prediction_reg[29]  ( .D(pc_out[29]), .CK(net19513), .RN(rst), 
        .Q(last_prediction[29]), .QN(n131) );
  DFFR_X1 \last_prediction_reg[6]  ( .D(pc_out[6]), .CK(net19518), .RN(rst), 
        .Q(last_prediction[6]), .QN(n129) );
  DFFS_X1 \last_prediction_reg[1]  ( .D(n585), .CK(net19518), .SN(rst), .Q(n85), .QN(last_prediction[1]) );
  DFFS_X1 \last_prediction_reg[0]  ( .D(n849), .CK(net19518), .SN(rst), .Q(n86), .QN(last_prediction[0]) );
  AND4_X1 U3 ( .A1(n165), .A2(n164), .A3(n167), .A4(n166), .ZN(n121) );
  OR2_X1 U4 ( .A1(n90), .A2(n108), .ZN(n194) );
  INV_X1 U5 ( .A(actual_addr[11]), .ZN(n272) );
  NAND2_X1 U6 ( .A1(actual_addr[18]), .A2(n77), .ZN(n76) );
  NAND2_X1 U7 ( .A1(actual_addr[17]), .A2(n79), .ZN(n78) );
  OAI22_X1 U8 ( .A1(n534), .A2(n382), .B1(n533), .B2(n468), .ZN(n9) );
  OAI21_X1 U9 ( .B1(n558), .B2(n526), .A(n9), .ZN(n10) );
  AOI222_X4 U10 ( .A1(n536), .A2(n553), .B1(n536), .B2(n10), .C1(n553), .C2(
        n10), .ZN(n380) );
  AOI21_X1 U11 ( .B1(n1475), .B2(n26), .A(n1474), .ZN(n11) );
  AOI22_X1 U12 ( .A1(n93), .A2(pc_in[5]), .B1(n249), .B2(n1480), .ZN(n12) );
  OAI211_X1 U13 ( .C1(n1481), .C2(n1584), .A(n11), .B(n12), .ZN(pc_out[5]) );
  NOR2_X1 U14 ( .A1(n884), .A2(n202), .ZN(n122) );
  AND2_X1 U15 ( .A1(n514), .A2(n552), .ZN(n13) );
  AOI211_X1 U16 ( .C1(n516), .C2(n515), .A(n13), .B(n513), .ZN(n14) );
  OAI211_X1 U17 ( .C1(n525), .C2(n521), .A(n520), .B(n519), .ZN(n15) );
  AOI21_X2 U18 ( .B1(n14), .B2(n15), .A(n522), .ZN(n592) );
  AOI22_X1 U19 ( .A1(actual_addr[20]), .A2(n74), .B1(n73), .B2(actual_addr[22]), .ZN(n70) );
  AOI22_X1 U20 ( .A1(n96), .A2(n1459), .B1(n93), .B2(pc_in[4]), .ZN(n16) );
  AOI21_X1 U21 ( .B1(n229), .B2(n1454), .A(n1453), .ZN(n17) );
  OAI211_X1 U22 ( .C1(n1460), .C2(n1584), .A(n16), .B(n17), .ZN(pc_out[4]) );
  NOR3_X1 U23 ( .A1(n884), .A2(n202), .A3(n807), .ZN(n141) );
  AOI211_X1 U24 ( .C1(n552), .C2(n553), .A(n550), .B(n551), .ZN(n18) );
  NAND3_X1 U25 ( .A1(n561), .A2(n562), .A3(n560), .ZN(n19) );
  AOI21_X1 U26 ( .B1(n18), .B2(n19), .A(n563), .ZN(n598) );
  NAND2_X1 U27 ( .A1(n606), .A2(n607), .ZN(N3360) );
  AOI22_X1 U28 ( .A1(n96), .A2(n1415), .B1(n93), .B2(pc_in[31]), .ZN(n20) );
  AOI21_X1 U29 ( .B1(n229), .B2(n1410), .A(n1409), .ZN(n21) );
  OAI211_X1 U30 ( .C1(n1416), .C2(n1584), .A(n20), .B(n21), .ZN(pc_out[31]) );
  AND4_X1 U31 ( .A1(n150), .A2(n147), .A3(n149), .A4(n148), .ZN(n22) );
  AND3_X1 U32 ( .A1(n896), .A2(n95), .A3(n900), .ZN(n1581) );
  INV_X1 U33 ( .A(n146), .ZN(n23) );
  INV_X1 U34 ( .A(misprediction_BAR), .ZN(n24) );
  AND3_X4 U35 ( .A1(n176), .A2(n175), .A3(n177), .ZN(n1584) );
  AOI22_X1 U36 ( .A1(n1371), .A2(n1370), .B1(n249), .B2(n1369), .ZN(n1372) );
  AND4_X2 U37 ( .A1(n152), .A2(n153), .A3(n151), .A4(n121), .ZN(n94) );
  NOR2_X1 U38 ( .A1(n886), .A2(n885), .ZN(n25) );
  NOR2_X1 U39 ( .A1(n886), .A2(n885), .ZN(n26) );
  CLKBUF_X3 U40 ( .A(n1567), .Z(n229) );
  AND3_X1 U41 ( .A1(n59), .A2(n1372), .A3(n28), .ZN(n27) );
  BUF_X2 U42 ( .A(n23), .Z(n201) );
  INV_X1 U43 ( .A(actual_addr[19]), .ZN(n281) );
  INV_X1 U44 ( .A(actual_addr[17]), .ZN(n278) );
  OR2_X1 U45 ( .A1(n247), .A2(pc_fetch[2]), .ZN(n28) );
  BUF_X4 U46 ( .A(n172), .Z(n93) );
  OR2_X1 U47 ( .A1(n1584), .A2(n1527), .ZN(n29) );
  OR2_X1 U48 ( .A1(n1584), .A2(n1439), .ZN(n30) );
  OR2_X1 U49 ( .A1(n1584), .A2(n1585), .ZN(n31) );
  OR2_X1 U50 ( .A1(n1584), .A2(n1550), .ZN(n32) );
  OR2_X1 U51 ( .A1(n1584), .A2(n1504), .ZN(n33) );
  INV_X1 U52 ( .A(actual_addr[18]), .ZN(n280) );
  INV_X4 U53 ( .A(n280), .ZN(n279) );
  OR2_X1 U54 ( .A1(n1350), .A2(n1584), .ZN(n61) );
  BUF_X1 U55 ( .A(n1581), .Z(n248) );
  BUF_X1 U56 ( .A(n1581), .Z(n96) );
  OR2_X1 U57 ( .A1(n1281), .A2(n1584), .ZN(n60) );
  INV_X1 U58 ( .A(n146), .ZN(n34) );
  INV_X2 U59 ( .A(n277), .ZN(n35) );
  CLKBUF_X3 U60 ( .A(n240), .Z(n239) );
  CLKBUF_X3 U61 ( .A(n244), .Z(n243) );
  CLKBUF_X2 U62 ( .A(n240), .Z(n55) );
  CLKBUF_X2 U63 ( .A(n244), .Z(n56) );
  CLKBUF_X3 U64 ( .A(n1569), .Z(n57) );
  BUF_X4 U65 ( .A(n1568), .Z(n36) );
  BUF_X4 U66 ( .A(n1570), .Z(n37) );
  BUF_X4 U67 ( .A(n1572), .Z(n38) );
  BUF_X4 U68 ( .A(n1574), .Z(n39) );
  BUF_X8 U69 ( .A(n1575), .Z(n40) );
  CLKBUF_X3 U70 ( .A(rst), .Z(n41) );
  INV_X2 U71 ( .A(n284), .ZN(n42) );
  INV_X2 U72 ( .A(n272), .ZN(n43) );
  INV_X2 U73 ( .A(n285), .ZN(n44) );
  INV_X2 U74 ( .A(n278), .ZN(n45) );
  INV_X2 U75 ( .A(n282), .ZN(n46) );
  INV_X2 U76 ( .A(n281), .ZN(n47) );
  INV_X2 U77 ( .A(n283), .ZN(n48) );
  INV_X2 U78 ( .A(n273), .ZN(n49) );
  INV_X2 U79 ( .A(n275), .ZN(n50) );
  INV_X2 U80 ( .A(n274), .ZN(n51) );
  INV_X1 U81 ( .A(actual_addr[16]), .ZN(n277) );
  INV_X2 U82 ( .A(n276), .ZN(n52) );
  NAND2_X1 U83 ( .A1(actual_addr[16]), .A2(n117), .ZN(n158) );
  NAND2_X1 U84 ( .A1(n367), .A2(n366), .ZN(n510) );
  BUF_X1 U85 ( .A(n57), .Z(n236) );
  BUF_X1 U86 ( .A(n57), .Z(n234) );
  INV_X1 U87 ( .A(actual_addr[22]), .ZN(n284) );
  INV_X1 U88 ( .A(actual_addr[20]), .ZN(n282) );
  NAND2_X1 U89 ( .A1(n877), .A2(last_prediction[0]), .ZN(n82) );
  OR2_X1 U90 ( .A1(n285), .A2(last_prediction[23]), .ZN(n155) );
  NAND2_X1 U91 ( .A1(n1120), .A2(last_prediction[1]), .ZN(n83) );
  OR2_X1 U92 ( .A1(n283), .A2(last_prediction[21]), .ZN(n154) );
  INV_X1 U93 ( .A(actual_addr[21]), .ZN(n283) );
  INV_X1 U94 ( .A(actual_addr[1]), .ZN(n1120) );
  INV_X1 U95 ( .A(actual_addr[23]), .ZN(n285) );
  INV_X1 U96 ( .A(actual_addr[15]), .ZN(n276) );
  INV_X1 U97 ( .A(actual_addr[13]), .ZN(n274) );
  INV_X1 U98 ( .A(actual_addr[14]), .ZN(n275) );
  INV_X1 U99 ( .A(actual_addr[12]), .ZN(n273) );
  OR2_X1 U100 ( .A1(n543), .A2(n544), .ZN(n540) );
  OR2_X1 U101 ( .A1(n564), .A2(n566), .ZN(n563) );
  OR2_X1 U102 ( .A1(n523), .A2(n524), .ZN(n522) );
  AND2_X1 U103 ( .A1(n538), .A2(n458), .ZN(n524) );
  AOI21_X1 U104 ( .B1(n375), .B2(\last_hit_index[2] ), .A(n474), .ZN(n482) );
  AND2_X1 U105 ( .A1(n538), .A2(n462), .ZN(n566) );
  INV_X1 U106 ( .A(n510), .ZN(n375) );
  AND2_X1 U107 ( .A1(n886), .A2(n200), .ZN(n81) );
  INV_X1 U108 ( .A(n901), .ZN(n95) );
  INV_X1 U109 ( .A(n607), .ZN(n587) );
  AOI21_X1 U110 ( .B1(n558), .B2(n556), .A(n550), .ZN(n446) );
  AND2_X1 U111 ( .A1(n370), .A2(n368), .ZN(n434) );
  INV_X1 U112 ( .A(n384), .ZN(n550) );
  INV_X1 U113 ( .A(n533), .ZN(n528) );
  INV_X1 U114 ( .A(n531), .ZN(n536) );
  INV_X1 U115 ( .A(n534), .ZN(n526) );
  INV_X1 U116 ( .A(n471), .ZN(n467) );
  INV_X1 U117 ( .A(n455), .ZN(n477) );
  NAND4_X1 U118 ( .A1(n342), .A2(n341), .A3(n340), .A4(n339), .ZN(n518) );
  NAND4_X1 U119 ( .A1(n309), .A2(n308), .A3(n307), .A4(n306), .ZN(n471) );
  NAND4_X1 U120 ( .A1(n346), .A2(n345), .A3(n344), .A4(n343), .ZN(n517) );
  NAND4_X1 U121 ( .A1(n333), .A2(n332), .A3(n331), .A4(n330), .ZN(n533) );
  INV_X1 U122 ( .A(n202), .ZN(n200) );
  BUF_X2 U123 ( .A(n1571), .Z(n240) );
  BUF_X2 U124 ( .A(n1573), .Z(n244) );
  BUF_X1 U125 ( .A(n1574), .Z(n246) );
  BUF_X1 U126 ( .A(n1568), .Z(n232) );
  INV_X1 U127 ( .A(n561), .ZN(n538) );
  INV_X1 U128 ( .A(n602), .ZN(n588) );
  INV_X1 U129 ( .A(n570), .ZN(n568) );
  INV_X1 U130 ( .A(n579), .ZN(n577) );
  INV_X1 U131 ( .A(n582), .ZN(n580) );
  NOR2_X2 U132 ( .A1(\last_set[1] ), .A2(n305), .ZN(n571) );
  INV_X1 U133 ( .A(n576), .ZN(n574) );
  INV_X1 U134 ( .A(n586), .ZN(n583) );
  NAND2_X1 U135 ( .A1(n508), .A2(\last_hit_index[2] ), .ZN(n561) );
  INV_X1 U136 ( .A(pc_fetch[10]), .ZN(n65) );
  NOR2_X1 U137 ( .A1(n109), .A2(n120), .ZN(n508) );
  INV_X1 U138 ( .A(pc_fetch[8]), .ZN(n66) );
  BUF_X1 U139 ( .A(n1), .Z(n257) );
  BUF_X1 U140 ( .A(n8), .Z(n250) );
  BUF_X1 U141 ( .A(n4), .Z(n254) );
  INV_X1 U142 ( .A(pc_fetch[3]), .ZN(n1586) );
  BUF_X1 U143 ( .A(n2), .Z(n256) );
  BUF_X1 U144 ( .A(n5), .Z(n253) );
  BUF_X1 U145 ( .A(n3), .Z(n255) );
  BUF_X1 U146 ( .A(n7), .Z(n251) );
  BUF_X1 U147 ( .A(n6), .Z(n252) );
  NAND3_X1 U148 ( .A1(n1502), .A2(n1503), .A3(n33), .ZN(pc_out[6]) );
  NAND3_X1 U149 ( .A1(n1548), .A2(n1549), .A3(n32), .ZN(pc_out[8]) );
  NAND3_X1 U150 ( .A1(n1582), .A2(n1583), .A3(n31), .ZN(pc_out[9]) );
  NAND3_X1 U151 ( .A1(n1438), .A2(n1437), .A3(n30), .ZN(pc_out[3]) );
  NAND3_X1 U152 ( .A1(n1526), .A2(n1525), .A3(n29), .ZN(pc_out[7]) );
  NOR2_X1 U153 ( .A1(n1226), .A2(n58), .ZN(n1234) );
  AND2_X1 U154 ( .A1(n1227), .A2(n26), .ZN(n58) );
  NAND3_X1 U155 ( .A1(n59), .A2(n1372), .A3(n28), .ZN(pc_out[2]) );
  INV_X1 U156 ( .A(n143), .ZN(n59) );
  NAND3_X1 U157 ( .A1(n1279), .A2(n1280), .A3(n60), .ZN(pc_out[26]) );
  NAND3_X1 U158 ( .A1(n1348), .A2(n1349), .A3(n61), .ZN(pc_out[29]) );
  NOR2_X1 U159 ( .A1(n1318), .A2(n62), .ZN(n1326) );
  AND2_X1 U160 ( .A1(n26), .A2(n1319), .ZN(n62) );
  NOR2_X1 U161 ( .A1(n1386), .A2(n63), .ZN(n1394) );
  AND2_X1 U162 ( .A1(n26), .A2(n1387), .ZN(n63) );
  NOR2_X1 U163 ( .A1(n1249), .A2(n68), .ZN(n1257) );
  AND2_X1 U164 ( .A1(n26), .A2(n1250), .ZN(n68) );
  NOR2_X1 U165 ( .A1(n1295), .A2(n69), .ZN(n1303) );
  AND2_X1 U166 ( .A1(n26), .A2(n1296), .ZN(n69) );
  NAND3_X1 U167 ( .A1(n155), .A2(n154), .A3(n70), .ZN(n89) );
  AOI22_X1 U168 ( .A1(actual_addr[0]), .A2(n86), .B1(actual_addr[1]), .B2(n85), 
        .ZN(n84) );
  NOR2_X1 U169 ( .A1(n72), .A2(n157), .ZN(n152) );
  NAND4_X1 U170 ( .A1(n76), .A2(n78), .A3(n158), .A4(n71), .ZN(n157) );
  NAND2_X1 U171 ( .A1(actual_addr[19]), .A2(n75), .ZN(n71) );
  NAND3_X1 U172 ( .A1(n154), .A2(n155), .A3(n70), .ZN(n72) );
  INV_X1 U173 ( .A(actual_addr[0]), .ZN(n877) );
  NAND2_X1 U174 ( .A1(n80), .A2(n197), .ZN(n896) );
  NAND3_X1 U175 ( .A1(n94), .A2(n90), .A3(n81), .ZN(n80) );
  NAND3_X1 U176 ( .A1(n82), .A2(n83), .A3(n84), .ZN(n502) );
  CLKBUF_X3 U177 ( .A(n303), .Z(n87) );
  CLKBUF_X3 U178 ( .A(n303), .Z(n88) );
  INV_X1 U179 ( .A(n34), .ZN(n303) );
  AND4_X1 U180 ( .A1(n150), .A2(n149), .A3(n148), .A4(n147), .ZN(n90) );
  INV_X1 U181 ( .A(n247), .ZN(n91) );
  NOR2_X1 U182 ( .A1(n157), .A2(n89), .ZN(n92) );
  INV_X1 U183 ( .A(n23), .ZN(misprediction_BAR) );
  INV_X1 U184 ( .A(n172), .ZN(n247) );
  CLKBUF_X3 U185 ( .A(n1567), .Z(n230) );
  CLKBUF_X3 U186 ( .A(n1581), .Z(n249) );
  BUF_X1 U187 ( .A(n590), .Z(n97) );
  BUF_X1 U188 ( .A(n590), .Z(n98) );
  AOI21_X1 U189 ( .B1(n171), .B2(n508), .A(n170), .ZN(n590) );
  BUF_X1 U190 ( .A(n599), .Z(n99) );
  BUF_X1 U191 ( .A(n599), .Z(n100) );
  AOI21_X1 U192 ( .B1(n171), .B2(n564), .A(n566), .ZN(n599) );
  BUF_X1 U193 ( .A(n593), .Z(n101) );
  BUF_X1 U194 ( .A(n593), .Z(n102) );
  AOI21_X1 U195 ( .B1(n171), .B2(n523), .A(n524), .ZN(n593) );
  BUF_X1 U196 ( .A(n596), .Z(n103) );
  BUF_X1 U197 ( .A(n596), .Z(n104) );
  AND2_X1 U198 ( .A1(n561), .A2(n34), .ZN(n171) );
  BUF_X2 U199 ( .A(rst), .Z(n304) );
  INV_X2 U200 ( .A(n271), .ZN(n270) );
  NAND2_X1 U201 ( .A1(n587), .A2(n566), .ZN(n601) );
  AOI21_X1 U202 ( .B1(n484), .B2(n483), .A(n482), .ZN(n589) );
  NAND2_X1 U203 ( .A1(n587), .A2(n524), .ZN(n594) );
  AOI21_X1 U204 ( .B1(n542), .B2(n541), .A(n540), .ZN(n595) );
  NAND2_X1 U205 ( .A1(n587), .A2(n544), .ZN(n597) );
  BUF_X2 U206 ( .A(n38), .Z(n241) );
  BUF_X2 U207 ( .A(n37), .Z(n237) );
  BUF_X2 U208 ( .A(n57), .Z(n233) );
  BUF_X2 U209 ( .A(n39), .Z(n245) );
  BUF_X2 U210 ( .A(n36), .Z(n231) );
  BUF_X2 U211 ( .A(n57), .Z(n235) );
  NOR2_X1 U212 ( .A1(n886), .A2(n885), .ZN(n1567) );
  AOI21_X1 U213 ( .B1(n171), .B2(n543), .A(n544), .ZN(n596) );
  NOR2_X1 U214 ( .A1(n561), .A2(n460), .ZN(n544) );
  OAI21_X1 U215 ( .B1(n355), .B2(n518), .A(n349), .ZN(n350) );
  OAI21_X1 U216 ( .B1(n380), .B2(n556), .A(n347), .ZN(n356) );
  OAI21_X1 U217 ( .B1(n380), .B2(n558), .A(n338), .ZN(n355) );
  INV_X1 U218 ( .A(n556), .ZN(n468) );
  INV_X1 U219 ( .A(n558), .ZN(n382) );
  NAND4_X1 U220 ( .A1(n329), .A2(n328), .A3(n327), .A4(n326), .ZN(n534) );
  NAND4_X1 U221 ( .A1(n325), .A2(n324), .A3(n323), .A4(n322), .ZN(n558) );
  NAND3_X1 U222 ( .A1(n106), .A2(\last_set[0] ), .A3(\last_set[1] ), .ZN(n579)
         );
  NAND2_X1 U223 ( .A1(\last_set[0] ), .A2(\last_set[2] ), .ZN(n305) );
  INV_X1 U224 ( .A(actual_addr[4]), .ZN(n261) );
  INV_X1 U225 ( .A(actual_addr[24]), .ZN(n287) );
  INV_X1 U226 ( .A(actual_addr[10]), .ZN(n271) );
  INV_X1 U227 ( .A(actual_addr[26]), .ZN(n291) );
  OR2_X1 U228 ( .A1(n276), .A2(last_prediction[15]), .ZN(n166) );
  OR2_X1 U229 ( .A1(n274), .A2(last_prediction[13]), .ZN(n167) );
  OR2_X1 U230 ( .A1(n275), .A2(last_prediction[14]), .ZN(n164) );
  OR2_X1 U231 ( .A1(n273), .A2(last_prediction[12]), .ZN(n165) );
  NOR2_X2 U232 ( .A1(n105), .A2(n305), .ZN(n509) );
  NAND3_X1 U233 ( .A1(n119), .A2(n106), .A3(\last_set[1] ), .ZN(n582) );
  NOR3_X1 U234 ( .A1(n381), .A2(n380), .A3(n510), .ZN(n462) );
  NAND4_X1 U235 ( .A1(n317), .A2(n316), .A3(n315), .A4(n314), .ZN(n553) );
  NAND4_X1 U236 ( .A1(n313), .A2(n312), .A3(n311), .A4(n310), .ZN(n531) );
  NAND3_X1 U237 ( .A1(n119), .A2(\last_set[1] ), .A3(\last_set[2] ), .ZN(n570)
         );
  BUF_X1 U238 ( .A(n1572), .Z(n242) );
  BUF_X1 U239 ( .A(n1570), .Z(n238) );
  NAND3_X1 U240 ( .A1(n105), .A2(n106), .A3(\last_set[0] ), .ZN(n586) );
  INV_X1 U241 ( .A(pc_fetch[4]), .ZN(n608) );
  NAND4_X1 U242 ( .A1(n321), .A2(n320), .A3(n319), .A4(n318), .ZN(n514) );
  NOR3_X1 U243 ( .A1(pc_fetch[4]), .A2(n1586), .A3(n609), .ZN(n1572) );
  NOR3_X1 U244 ( .A1(pc_fetch[2]), .A2(pc_fetch[4]), .A3(n1586), .ZN(n1573) );
  NOR3_X1 U245 ( .A1(pc_fetch[3]), .A2(n609), .A3(n608), .ZN(n1570) );
  NOR3_X1 U246 ( .A1(pc_fetch[2]), .A2(pc_fetch[3]), .A3(n608), .ZN(n1571) );
  INV_X1 U247 ( .A(pc_fetch[2]), .ZN(n609) );
  INV_X1 U248 ( .A(n514), .ZN(n516) );
  INV_X1 U249 ( .A(n370), .ZN(n480) );
  NOR2_X1 U250 ( .A1(n531), .A2(n553), .ZN(n364) );
  NAND2_X1 U251 ( .A1(verify), .A2(ID_EN), .ZN(n607) );
  NAND4_X1 U252 ( .A1(n363), .A2(n362), .A3(n361), .A4(n360), .ZN(n465) );
  INV_X2 U253 ( .A(n258), .ZN(n212) );
  INV_X2 U254 ( .A(n259), .ZN(n216) );
  INV_X2 U255 ( .A(n261), .ZN(n260) );
  INV_X2 U256 ( .A(n268), .ZN(n222) );
  INV_X2 U257 ( .A(n263), .ZN(n262) );
  INV_X2 U258 ( .A(n265), .ZN(n264) );
  INV_X2 U259 ( .A(n267), .ZN(n266) );
  INV_X2 U260 ( .A(n269), .ZN(n204) );
  INV_X2 U261 ( .A(n301), .ZN(n300) );
  BUF_X2 U262 ( .A(n1563), .Z(n228) );
  INV_X2 U263 ( .A(n299), .ZN(n298) );
  INV_X2 U264 ( .A(n297), .ZN(n296) );
  INV_X2 U265 ( .A(n295), .ZN(n294) );
  INV_X2 U266 ( .A(n293), .ZN(n292) );
  INV_X2 U267 ( .A(n291), .ZN(n290) );
  INV_X2 U268 ( .A(n289), .ZN(n288) );
  INV_X2 U269 ( .A(n287), .ZN(n286) );
  BUF_X2 U270 ( .A(n1563), .Z(n227) );
  BUF_X2 U271 ( .A(n1563), .Z(n226) );
  NAND4_X2 U272 ( .A1(n337), .A2(n336), .A3(n335), .A4(n334), .ZN(n556) );
  NOR2_X1 U273 ( .A1(\last_hit_index[0] ), .A2(\last_hit_index[1] ), .ZN(n564)
         );
  NOR2_X1 U274 ( .A1(\last_hit_index[1] ), .A2(n109), .ZN(n543) );
  NOR2_X1 U275 ( .A1(\last_hit_index[0] ), .A2(n120), .ZN(n523) );
  NAND2_X1 U276 ( .A1(n196), .A2(n199), .ZN(n882) );
  NAND2_X1 U277 ( .A1(n201), .A2(n212), .ZN(n211) );
  OAI21_X1 U278 ( .B1(n228), .B2(n1429), .A(n215), .ZN(n1430) );
  NAND2_X1 U279 ( .A1(n201), .A2(n216), .ZN(n215) );
  OAI21_X1 U280 ( .B1(n227), .B2(n1452), .A(n217), .ZN(n1453) );
  NAND2_X1 U281 ( .A1(n201), .A2(n260), .ZN(n217) );
  OAI21_X1 U282 ( .B1(n228), .B2(n1540), .A(n221), .ZN(n1541) );
  NAND2_X1 U283 ( .A1(n201), .A2(n222), .ZN(n221) );
  OAI21_X1 U284 ( .B1(n227), .B2(n1473), .A(n218), .ZN(n1474) );
  NAND2_X1 U285 ( .A1(n201), .A2(n262), .ZN(n218) );
  OAI21_X1 U286 ( .B1(n228), .B2(n1494), .A(n219), .ZN(n1495) );
  NAND2_X1 U287 ( .A1(n201), .A2(n264), .ZN(n219) );
  OAI21_X1 U288 ( .B1(n227), .B2(n1517), .A(n220), .ZN(n1518) );
  NAND2_X1 U289 ( .A1(n201), .A2(n266), .ZN(n220) );
  OAI21_X1 U290 ( .B1(n228), .B2(n1564), .A(n203), .ZN(n1565) );
  NAND2_X1 U291 ( .A1(n201), .A2(n204), .ZN(n203) );
  NOR2_X1 U292 ( .A1(n375), .A2(n561), .ZN(n170) );
  OAI21_X1 U293 ( .B1(n227), .B2(n1408), .A(n214), .ZN(n1409) );
  NAND2_X1 U294 ( .A1(n201), .A2(n300), .ZN(n214) );
  OAI21_X1 U295 ( .B1(n227), .B2(n1385), .A(n213), .ZN(n1386) );
  NAND2_X1 U296 ( .A1(n24), .A2(n298), .ZN(n213) );
  OAI21_X1 U297 ( .B1(n228), .B2(n1340), .A(n210), .ZN(n1341) );
  NAND2_X1 U298 ( .A1(n201), .A2(n296), .ZN(n210) );
  OAI21_X1 U299 ( .B1(n227), .B2(n1317), .A(n209), .ZN(n1318) );
  NAND2_X1 U300 ( .A1(n24), .A2(n294), .ZN(n209) );
  OAI21_X1 U301 ( .B1(n228), .B2(n1294), .A(n208), .ZN(n1295) );
  NAND2_X1 U302 ( .A1(n24), .A2(n292), .ZN(n208) );
  OAI21_X1 U303 ( .B1(n227), .B2(n1271), .A(n207), .ZN(n1272) );
  NAND2_X1 U304 ( .A1(n201), .A2(n290), .ZN(n207) );
  OAI21_X1 U305 ( .B1(n228), .B2(n1248), .A(n206), .ZN(n1249) );
  NAND2_X1 U306 ( .A1(n24), .A2(n288), .ZN(n206) );
  OAI21_X1 U307 ( .B1(n228), .B2(n1225), .A(n205), .ZN(n1226) );
  NAND2_X1 U308 ( .A1(n24), .A2(n286), .ZN(n205) );
  OAI21_X1 U309 ( .B1(n23), .B2(n906), .A(n173), .ZN(n172) );
  NAND4_X1 U310 ( .A1(n195), .A2(n194), .A3(n200), .A4(n193), .ZN(n173) );
  OR2_X1 U311 ( .A1(n94), .A2(n108), .ZN(n195) );
  INV_X1 U312 ( .A(n199), .ZN(n198) );
  NAND2_X1 U313 ( .A1(n108), .A2(n200), .ZN(n199) );
  INV_X1 U314 ( .A(n883), .ZN(n193) );
  OAI22_X1 U315 ( .A1(actual_addr[5]), .A2(n115), .B1(actual_addr[4]), .B2(
        n136), .ZN(n169) );
  OAI22_X1 U316 ( .A1(actual_addr[25]), .A2(n116), .B1(actual_addr[24]), .B2(
        n137), .ZN(n174) );
  OAI22_X1 U317 ( .A1(actual_addr[11]), .A2(n114), .B1(actual_addr[10]), .B2(
        n135), .ZN(n168) );
  NOR2_X1 U318 ( .A1(n190), .A2(n189), .ZN(n490) );
  NOR2_X1 U319 ( .A1(actual_addr[26]), .A2(n130), .ZN(n189) );
  NOR2_X1 U320 ( .A1(actual_addr[27]), .A2(n134), .ZN(n190) );
  NOR2_X1 U321 ( .A1(n183), .A2(n182), .ZN(n491) );
  NOR2_X1 U322 ( .A1(actual_addr[28]), .A2(n127), .ZN(n182) );
  NOR2_X1 U323 ( .A1(actual_addr[29]), .A2(n131), .ZN(n183) );
  NOR2_X1 U324 ( .A1(n186), .A2(n187), .ZN(n499) );
  NOR2_X1 U325 ( .A1(actual_addr[6]), .A2(n129), .ZN(n186) );
  NOR2_X1 U326 ( .A1(actual_addr[7]), .A2(n133), .ZN(n187) );
  NOR2_X1 U327 ( .A1(n185), .A2(n184), .ZN(n492) );
  NOR2_X1 U328 ( .A1(actual_addr[30]), .A2(n128), .ZN(n184) );
  NOR2_X1 U329 ( .A1(actual_addr[31]), .A2(n132), .ZN(n185) );
  INV_X1 U330 ( .A(n179), .ZN(n504) );
  OAI22_X1 U331 ( .A1(actual_addr[12]), .A2(n112), .B1(actual_addr[13]), .B2(
        n125), .ZN(n179) );
  INV_X1 U332 ( .A(n178), .ZN(n485) );
  OAI22_X1 U333 ( .A1(actual_addr[16]), .A2(n117), .B1(actual_addr[17]), .B2(
        n79), .ZN(n178) );
  INV_X1 U334 ( .A(n181), .ZN(n505) );
  OAI22_X1 U335 ( .A1(actual_addr[14]), .A2(n113), .B1(actual_addr[15]), .B2(
        n126), .ZN(n181) );
  INV_X1 U336 ( .A(n180), .ZN(n486) );
  OAI22_X1 U337 ( .A1(actual_addr[18]), .A2(n77), .B1(actual_addr[19]), .B2(
        n75), .ZN(n180) );
  NAND2_X1 U338 ( .A1(n145), .A2(n144), .ZN(n156) );
  AOI22_X1 U339 ( .A1(actual_addr[2]), .A2(n110), .B1(actual_addr[8]), .B2(
        n123), .ZN(n144) );
  AOI22_X1 U340 ( .A1(actual_addr[3]), .A2(n111), .B1(actual_addr[9]), .B2(
        n124), .ZN(n145) );
  NOR2_X1 U341 ( .A1(n192), .A2(n191), .ZN(n487) );
  NOR2_X1 U342 ( .A1(actual_addr[20]), .A2(n74), .ZN(n191) );
  NOR2_X1 U343 ( .A1(actual_addr[21]), .A2(n138), .ZN(n192) );
  INV_X1 U344 ( .A(n223), .ZN(n507) );
  OAI22_X1 U345 ( .A1(actual_addr[8]), .A2(n123), .B1(actual_addr[9]), .B2(
        n124), .ZN(n223) );
  INV_X1 U346 ( .A(n188), .ZN(n506) );
  OAI22_X1 U347 ( .A1(actual_addr[2]), .A2(n110), .B1(actual_addr[3]), .B2(
        n111), .ZN(n188) );
  NOR2_X1 U348 ( .A1(n225), .A2(n224), .ZN(n488) );
  NOR2_X1 U349 ( .A1(actual_addr[22]), .A2(n73), .ZN(n224) );
  NOR2_X1 U350 ( .A1(actual_addr[23]), .A2(n139), .ZN(n225) );
  AND2_X1 U351 ( .A1(n193), .A2(n122), .ZN(n107) );
  NOR2_X1 U352 ( .A1(n197), .A2(n884), .ZN(n118) );
  INV_X1 U353 ( .A(actual_addr[3]), .ZN(n259) );
  INV_X1 U354 ( .A(actual_addr[2]), .ZN(n258) );
  INV_X1 U355 ( .A(actual_addr[9]), .ZN(n269) );
  INV_X1 U356 ( .A(actual_addr[8]), .ZN(n268) );
  INV_X1 U357 ( .A(actual_addr[6]), .ZN(n265) );
  INV_X1 U358 ( .A(actual_addr[28]), .ZN(n295) );
  INV_X1 U359 ( .A(actual_addr[30]), .ZN(n299) );
  INV_X1 U360 ( .A(actual_addr[27]), .ZN(n293) );
  INV_X1 U361 ( .A(actual_addr[7]), .ZN(n267) );
  INV_X1 U362 ( .A(actual_addr[29]), .ZN(n297) );
  INV_X1 U363 ( .A(actual_addr[31]), .ZN(n301) );
  INV_X1 U364 ( .A(actual_addr[25]), .ZN(n289) );
  INV_X1 U365 ( .A(actual_addr[5]), .ZN(n263) );
  NAND2_X1 U366 ( .A1(n886), .A2(n198), .ZN(n197) );
  AND2_X1 U367 ( .A1(n122), .A2(n108), .ZN(n140) );
  OAI211_X1 U368 ( .C1(n1359), .C2(n227), .A(n142), .B(n211), .ZN(n143) );
  NAND2_X1 U369 ( .A1(n25), .A2(n1360), .ZN(n142) );
  OAI21_X1 U370 ( .B1(n160), .B2(n159), .A(verify), .ZN(n146) );
  NAND4_X1 U371 ( .A1(n92), .A2(n153), .A3(n151), .A4(n121), .ZN(n160) );
  NAND4_X1 U372 ( .A1(n150), .A2(n147), .A3(n149), .A4(n148), .ZN(n159) );
  NOR2_X1 U373 ( .A1(n502), .A2(n501), .ZN(n147) );
  NOR2_X1 U374 ( .A1(n503), .A2(n496), .ZN(n148) );
  NOR2_X1 U375 ( .A1(n494), .A2(n495), .ZN(n149) );
  NOR2_X1 U376 ( .A1(n493), .A2(n500), .ZN(n150) );
  NOR2_X1 U377 ( .A1(n161), .A2(n162), .ZN(n151) );
  NOR2_X1 U378 ( .A1(n163), .A2(n156), .ZN(n153) );
  NAND2_X1 U379 ( .A1(n486), .A2(n505), .ZN(n161) );
  NAND2_X1 U380 ( .A1(n485), .A2(n504), .ZN(n162) );
  NAND4_X1 U381 ( .A1(n488), .A2(n506), .A3(n507), .A4(n487), .ZN(n163) );
  INV_X1 U382 ( .A(n168), .ZN(n497) );
  INV_X1 U383 ( .A(n169), .ZN(n498) );
  INV_X1 U384 ( .A(n174), .ZN(n489) );
  NAND3_X1 U385 ( .A1(n94), .A2(n22), .A3(n141), .ZN(n175) );
  NAND3_X1 U386 ( .A1(n94), .A2(n22), .A3(n107), .ZN(n176) );
  AOI21_X1 U387 ( .B1(n193), .B2(n140), .A(n118), .ZN(n177) );
  INV_X1 U388 ( .A(n1584), .ZN(n1371) );
  NAND3_X1 U389 ( .A1(n195), .A2(n200), .A3(n194), .ZN(n885) );
  NAND3_X1 U390 ( .A1(n94), .A2(n22), .A3(n200), .ZN(n196) );
  INV_X1 U391 ( .A(n906), .ZN(n202) );
  NAND3_X1 U392 ( .A1(n105), .A2(n119), .A3(n106), .ZN(n602) );
  AOI22_X1 U393 ( .A1(n588), .A2(\cache[0][3][YOUTH][0] ), .B1(n509), .B2(
        \cache[7][3][YOUTH][0] ), .ZN(n309) );
  AOI22_X1 U394 ( .A1(n568), .A2(\cache[6][3][YOUTH][0] ), .B1(n577), .B2(
        \cache[3][3][YOUTH][0] ), .ZN(n308) );
  AOI22_X1 U395 ( .A1(n580), .A2(\cache[2][3][YOUTH][0] ), .B1(n571), .B2(
        \cache[5][3][YOUTH][0] ), .ZN(n307) );
  NAND3_X1 U396 ( .A1(n105), .A2(n119), .A3(\last_set[2] ), .ZN(n576) );
  AOI22_X1 U397 ( .A1(n574), .A2(\cache[4][3][YOUTH][0] ), .B1(n583), .B2(
        \cache[1][3][YOUTH][0] ), .ZN(n306) );
  AOI22_X1 U398 ( .A1(\cache[0][1][YOUTH][2] ), .A2(n588), .B1(
        \cache[7][1][YOUTH][2] ), .B2(n509), .ZN(n313) );
  AOI22_X1 U399 ( .A1(\cache[6][1][YOUTH][2] ), .A2(n568), .B1(
        \cache[3][1][YOUTH][2] ), .B2(n577), .ZN(n312) );
  AOI22_X1 U400 ( .A1(\cache[2][1][YOUTH][2] ), .A2(n580), .B1(
        \cache[5][1][YOUTH][2] ), .B2(n571), .ZN(n311) );
  AOI22_X1 U401 ( .A1(\cache[4][1][YOUTH][2] ), .A2(n574), .B1(
        \cache[1][1][YOUTH][2] ), .B2(n583), .ZN(n310) );
  AOI22_X1 U402 ( .A1(n588), .A2(\cache[0][0][YOUTH][2] ), .B1(n509), .B2(
        \cache[7][0][YOUTH][2] ), .ZN(n317) );
  AOI22_X1 U403 ( .A1(n568), .A2(\cache[6][0][YOUTH][2] ), .B1(n577), .B2(
        \cache[3][0][YOUTH][2] ), .ZN(n316) );
  AOI22_X1 U404 ( .A1(n580), .A2(\cache[2][0][YOUTH][2] ), .B1(n571), .B2(
        \cache[5][0][YOUTH][2] ), .ZN(n315) );
  AOI22_X1 U405 ( .A1(n574), .A2(\cache[4][0][YOUTH][2] ), .B1(n583), .B2(
        \cache[1][0][YOUTH][2] ), .ZN(n314) );
  AOI22_X1 U406 ( .A1(n588), .A2(\cache[0][2][YOUTH][2] ), .B1(n509), .B2(
        \cache[7][2][YOUTH][2] ), .ZN(n321) );
  AOI22_X1 U407 ( .A1(n568), .A2(\cache[6][2][YOUTH][2] ), .B1(n577), .B2(
        \cache[3][2][YOUTH][2] ), .ZN(n320) );
  AOI22_X1 U408 ( .A1(n580), .A2(\cache[2][2][YOUTH][2] ), .B1(n571), .B2(
        \cache[5][2][YOUTH][2] ), .ZN(n319) );
  AOI22_X1 U409 ( .A1(n574), .A2(\cache[4][2][YOUTH][2] ), .B1(n583), .B2(
        \cache[1][2][YOUTH][2] ), .ZN(n318) );
  AOI22_X1 U410 ( .A1(n588), .A2(\cache[0][0][YOUTH][1] ), .B1(n509), .B2(
        \cache[7][0][YOUTH][1] ), .ZN(n325) );
  AOI22_X1 U411 ( .A1(n568), .A2(\cache[6][0][YOUTH][1] ), .B1(n577), .B2(
        \cache[3][0][YOUTH][1] ), .ZN(n324) );
  AOI22_X1 U412 ( .A1(n580), .A2(\cache[2][0][YOUTH][1] ), .B1(n571), .B2(
        \cache[5][0][YOUTH][1] ), .ZN(n323) );
  AOI22_X1 U413 ( .A1(n574), .A2(\cache[4][0][YOUTH][1] ), .B1(n583), .B2(
        \cache[1][0][YOUTH][1] ), .ZN(n322) );
  AOI22_X1 U414 ( .A1(n588), .A2(\cache[0][1][YOUTH][1] ), .B1(n509), .B2(
        \cache[7][1][YOUTH][1] ), .ZN(n329) );
  AOI22_X1 U415 ( .A1(n568), .A2(\cache[6][1][YOUTH][1] ), .B1(n577), .B2(
        \cache[3][1][YOUTH][1] ), .ZN(n328) );
  AOI22_X1 U416 ( .A1(n580), .A2(\cache[2][1][YOUTH][1] ), .B1(n571), .B2(
        \cache[5][1][YOUTH][1] ), .ZN(n327) );
  AOI22_X1 U417 ( .A1(n574), .A2(\cache[4][1][YOUTH][1] ), .B1(n583), .B2(
        \cache[1][1][YOUTH][1] ), .ZN(n326) );
  AOI22_X1 U418 ( .A1(n588), .A2(\cache[0][1][YOUTH][0] ), .B1(n509), .B2(
        \cache[7][1][YOUTH][0] ), .ZN(n333) );
  AOI22_X1 U419 ( .A1(n568), .A2(\cache[6][1][YOUTH][0] ), .B1(n577), .B2(
        \cache[3][1][YOUTH][0] ), .ZN(n332) );
  AOI22_X1 U420 ( .A1(n580), .A2(\cache[2][1][YOUTH][0] ), .B1(n571), .B2(
        \cache[5][1][YOUTH][0] ), .ZN(n331) );
  AOI22_X1 U421 ( .A1(n574), .A2(\cache[4][1][YOUTH][0] ), .B1(n583), .B2(
        \cache[1][1][YOUTH][0] ), .ZN(n330) );
  AOI22_X1 U422 ( .A1(n588), .A2(\cache[0][0][YOUTH][0] ), .B1(n509), .B2(
        \cache[7][0][YOUTH][0] ), .ZN(n337) );
  AOI22_X1 U423 ( .A1(n568), .A2(\cache[6][0][YOUTH][0] ), .B1(n577), .B2(
        \cache[3][0][YOUTH][0] ), .ZN(n336) );
  AOI22_X1 U424 ( .A1(n580), .A2(\cache[2][0][YOUTH][0] ), .B1(n571), .B2(
        \cache[5][0][YOUTH][0] ), .ZN(n335) );
  AOI22_X1 U425 ( .A1(n574), .A2(\cache[4][0][YOUTH][0] ), .B1(n583), .B2(
        \cache[1][0][YOUTH][0] ), .ZN(n334) );
  NAND2_X1 U426 ( .A1(n380), .A2(n526), .ZN(n338) );
  AOI22_X1 U427 ( .A1(n588), .A2(\cache[0][2][YOUTH][1] ), .B1(n509), .B2(
        \cache[7][2][YOUTH][1] ), .ZN(n342) );
  AOI22_X1 U428 ( .A1(n568), .A2(\cache[6][2][YOUTH][1] ), .B1(n577), .B2(
        \cache[3][2][YOUTH][1] ), .ZN(n341) );
  AOI22_X1 U429 ( .A1(n580), .A2(\cache[2][2][YOUTH][1] ), .B1(n571), .B2(
        \cache[5][2][YOUTH][1] ), .ZN(n340) );
  AOI22_X1 U430 ( .A1(n574), .A2(\cache[4][2][YOUTH][1] ), .B1(n583), .B2(
        \cache[1][2][YOUTH][1] ), .ZN(n339) );
  AOI22_X1 U431 ( .A1(n588), .A2(\cache[0][2][YOUTH][0] ), .B1(n509), .B2(
        \cache[7][2][YOUTH][0] ), .ZN(n346) );
  AOI22_X1 U432 ( .A1(n568), .A2(\cache[6][2][YOUTH][0] ), .B1(n577), .B2(
        \cache[3][2][YOUTH][0] ), .ZN(n345) );
  AOI22_X1 U433 ( .A1(n580), .A2(\cache[2][2][YOUTH][0] ), .B1(n571), .B2(
        \cache[5][2][YOUTH][0] ), .ZN(n344) );
  AOI22_X1 U434 ( .A1(n574), .A2(\cache[4][2][YOUTH][0] ), .B1(n583), .B2(
        \cache[1][2][YOUTH][0] ), .ZN(n343) );
  NAND2_X1 U435 ( .A1(n380), .A2(n528), .ZN(n347) );
  AOI211_X1 U436 ( .C1(n518), .C2(n355), .A(n517), .B(n356), .ZN(n348) );
  INV_X1 U437 ( .A(n348), .ZN(n349) );
  AOI222_X1 U438 ( .A1(n364), .A2(n514), .B1(n364), .B2(n350), .C1(n514), .C2(
        n350), .ZN(n376) );
  INV_X1 U439 ( .A(n376), .ZN(n381) );
  AOI22_X1 U440 ( .A1(n588), .A2(\cache[0][3][YOUTH][1] ), .B1(n509), .B2(
        \cache[7][3][YOUTH][1] ), .ZN(n354) );
  AOI22_X1 U441 ( .A1(n568), .A2(\cache[6][3][YOUTH][1] ), .B1(n577), .B2(
        \cache[3][3][YOUTH][1] ), .ZN(n353) );
  AOI22_X1 U442 ( .A1(n580), .A2(\cache[2][3][YOUTH][1] ), .B1(n571), .B2(
        \cache[5][3][YOUTH][1] ), .ZN(n352) );
  AOI22_X1 U443 ( .A1(n574), .A2(\cache[4][3][YOUTH][1] ), .B1(n583), .B2(
        \cache[1][3][YOUTH][1] ), .ZN(n351) );
  NAND4_X1 U444 ( .A1(n354), .A2(n353), .A3(n352), .A4(n351), .ZN(n455) );
  NAND2_X1 U445 ( .A1(n477), .A2(n467), .ZN(n370) );
  AOI222_X1 U446 ( .A1(n518), .A2(n517), .B1(n518), .B2(n477), .C1(n517), .C2(
        n480), .ZN(n359) );
  AOI222_X1 U447 ( .A1(n356), .A2(n355), .B1(n356), .B2(n455), .C1(n355), .C2(
        n370), .ZN(n357) );
  NAND2_X1 U448 ( .A1(n455), .A2(n471), .ZN(n368) );
  OAI21_X1 U449 ( .B1(n357), .B2(n381), .A(n368), .ZN(n358) );
  AOI21_X1 U450 ( .B1(n381), .B2(n359), .A(n358), .ZN(n365) );
  AOI22_X1 U451 ( .A1(n588), .A2(\cache[0][3][YOUTH][2] ), .B1(n509), .B2(
        \cache[7][3][YOUTH][2] ), .ZN(n363) );
  AOI22_X1 U452 ( .A1(n568), .A2(\cache[6][3][YOUTH][2] ), .B1(n577), .B2(
        \cache[3][3][YOUTH][2] ), .ZN(n362) );
  AOI22_X1 U453 ( .A1(n580), .A2(\cache[2][3][YOUTH][2] ), .B1(n571), .B2(
        \cache[5][3][YOUTH][2] ), .ZN(n361) );
  AOI22_X1 U454 ( .A1(n574), .A2(\cache[4][3][YOUTH][2] ), .B1(n583), .B2(
        \cache[1][3][YOUTH][2] ), .ZN(n360) );
  OAI211_X1 U455 ( .C1(n365), .C2(n465), .A(n516), .B(n364), .ZN(n367) );
  NAND2_X1 U456 ( .A1(n365), .A2(n465), .ZN(n366) );
  INV_X1 U457 ( .A(n508), .ZN(n474) );
  NAND2_X1 U458 ( .A1(n509), .A2(n482), .ZN(n369) );
  NAND2_X1 U459 ( .A1(n471), .A2(n369), .ZN(N2805) );
  NAND2_X1 U460 ( .A1(n434), .A2(n369), .ZN(N2806) );
  INV_X1 U461 ( .A(n369), .ZN(n371) );
  INV_X1 U462 ( .A(n465), .ZN(n481) );
  AOI22_X1 U463 ( .A1(n480), .A2(n481), .B1(n465), .B2(n370), .ZN(n437) );
  NOR2_X1 U464 ( .A1(n371), .A2(n437), .ZN(N2807) );
  NOR2_X1 U465 ( .A1(n376), .A2(n510), .ZN(n458) );
  NAND2_X1 U466 ( .A1(n509), .A2(n522), .ZN(n372) );
  NAND2_X1 U467 ( .A1(n517), .A2(n372), .ZN(N2811) );
  NOR2_X1 U468 ( .A1(n518), .A2(n517), .ZN(n515) );
  AOI21_X1 U469 ( .B1(n518), .B2(n517), .A(n515), .ZN(n438) );
  NAND2_X1 U470 ( .A1(n438), .A2(n372), .ZN(N2812) );
  INV_X1 U471 ( .A(n372), .ZN(n374) );
  INV_X1 U472 ( .A(n515), .ZN(n373) );
  AOI22_X1 U473 ( .A1(n516), .A2(n515), .B1(n373), .B2(n514), .ZN(n441) );
  NOR2_X1 U474 ( .A1(n374), .A2(n441), .ZN(N2813) );
  NAND3_X1 U475 ( .A1(n380), .A2(n376), .A3(n375), .ZN(n460) );
  NAND2_X1 U476 ( .A1(n509), .A2(n540), .ZN(n377) );
  NAND2_X1 U477 ( .A1(n533), .A2(n377), .ZN(N2817) );
  NAND2_X1 U478 ( .A1(n526), .A2(n528), .ZN(n378) );
  INV_X1 U479 ( .A(n378), .ZN(n532) );
  AOI21_X1 U480 ( .B1(n534), .B2(n533), .A(n532), .ZN(n442) );
  NAND2_X1 U481 ( .A1(n442), .A2(n377), .ZN(N2818) );
  INV_X1 U482 ( .A(n377), .ZN(n379) );
  AOI22_X1 U483 ( .A1(n536), .A2(n532), .B1(n378), .B2(n531), .ZN(n445) );
  NOR2_X1 U484 ( .A1(n379), .A2(n445), .ZN(N2819) );
  NAND2_X1 U485 ( .A1(n509), .A2(n563), .ZN(n383) );
  NAND2_X1 U486 ( .A1(n556), .A2(n383), .ZN(N2823) );
  NAND2_X1 U487 ( .A1(n382), .A2(n468), .ZN(n384) );
  NAND2_X1 U488 ( .A1(n446), .A2(n383), .ZN(N2824) );
  INV_X1 U489 ( .A(n383), .ZN(n385) );
  INV_X1 U490 ( .A(n553), .ZN(n555) );
  AOI22_X1 U491 ( .A1(n555), .A2(n550), .B1(n384), .B2(n553), .ZN(n449) );
  NOR2_X1 U492 ( .A1(n385), .A2(n449), .ZN(N2825) );
  NAND2_X1 U493 ( .A1(n568), .A2(n482), .ZN(n386) );
  NAND2_X1 U494 ( .A1(n471), .A2(n386), .ZN(N2829) );
  NAND2_X1 U495 ( .A1(n434), .A2(n386), .ZN(N2830) );
  INV_X1 U496 ( .A(n386), .ZN(n387) );
  NOR2_X1 U497 ( .A1(n437), .A2(n387), .ZN(N2831) );
  NAND2_X1 U498 ( .A1(n568), .A2(n522), .ZN(n388) );
  NAND2_X1 U499 ( .A1(n517), .A2(n388), .ZN(N2835) );
  NAND2_X1 U500 ( .A1(n438), .A2(n388), .ZN(N2836) );
  INV_X1 U501 ( .A(n388), .ZN(n389) );
  NOR2_X1 U502 ( .A1(n441), .A2(n389), .ZN(N2837) );
  NAND2_X1 U503 ( .A1(n568), .A2(n540), .ZN(n390) );
  NAND2_X1 U504 ( .A1(n533), .A2(n390), .ZN(N2841) );
  NAND2_X1 U505 ( .A1(n442), .A2(n390), .ZN(N2842) );
  INV_X1 U506 ( .A(n390), .ZN(n391) );
  NOR2_X1 U507 ( .A1(n445), .A2(n391), .ZN(N2843) );
  NAND2_X1 U508 ( .A1(n568), .A2(n563), .ZN(n392) );
  NAND2_X1 U509 ( .A1(n556), .A2(n392), .ZN(N2847) );
  NAND2_X1 U510 ( .A1(n446), .A2(n392), .ZN(N2848) );
  INV_X1 U511 ( .A(n392), .ZN(n393) );
  NOR2_X1 U512 ( .A1(n449), .A2(n393), .ZN(N2849) );
  NAND2_X1 U513 ( .A1(n571), .A2(n482), .ZN(n394) );
  NAND2_X1 U514 ( .A1(n471), .A2(n394), .ZN(N2853) );
  NAND2_X1 U515 ( .A1(n434), .A2(n394), .ZN(N2854) );
  INV_X1 U516 ( .A(n394), .ZN(n395) );
  NOR2_X1 U517 ( .A1(n437), .A2(n395), .ZN(N2855) );
  NAND2_X1 U518 ( .A1(n571), .A2(n522), .ZN(n396) );
  NAND2_X1 U519 ( .A1(n517), .A2(n396), .ZN(N2859) );
  NAND2_X1 U520 ( .A1(n438), .A2(n396), .ZN(N2860) );
  INV_X1 U521 ( .A(n396), .ZN(n397) );
  NOR2_X1 U522 ( .A1(n441), .A2(n397), .ZN(N2861) );
  NAND2_X1 U523 ( .A1(n571), .A2(n540), .ZN(n398) );
  NAND2_X1 U524 ( .A1(n533), .A2(n398), .ZN(N2865) );
  NAND2_X1 U525 ( .A1(n442), .A2(n398), .ZN(N2866) );
  INV_X1 U526 ( .A(n398), .ZN(n399) );
  NOR2_X1 U527 ( .A1(n445), .A2(n399), .ZN(N2867) );
  NAND2_X1 U528 ( .A1(n571), .A2(n563), .ZN(n400) );
  NAND2_X1 U529 ( .A1(n556), .A2(n400), .ZN(N2871) );
  NAND2_X1 U530 ( .A1(n446), .A2(n400), .ZN(N2872) );
  INV_X1 U531 ( .A(n400), .ZN(n401) );
  NOR2_X1 U532 ( .A1(n449), .A2(n401), .ZN(N2873) );
  NAND2_X1 U533 ( .A1(n574), .A2(n482), .ZN(n402) );
  NAND2_X1 U534 ( .A1(n471), .A2(n402), .ZN(N2877) );
  NAND2_X1 U535 ( .A1(n434), .A2(n402), .ZN(N2878) );
  INV_X1 U536 ( .A(n402), .ZN(n403) );
  NOR2_X1 U537 ( .A1(n437), .A2(n403), .ZN(N2879) );
  NAND2_X1 U538 ( .A1(n574), .A2(n522), .ZN(n404) );
  NAND2_X1 U539 ( .A1(n517), .A2(n404), .ZN(N2883) );
  NAND2_X1 U540 ( .A1(n438), .A2(n404), .ZN(N2884) );
  INV_X1 U541 ( .A(n404), .ZN(n405) );
  NOR2_X1 U542 ( .A1(n441), .A2(n405), .ZN(N2885) );
  NAND2_X1 U543 ( .A1(n574), .A2(n540), .ZN(n406) );
  NAND2_X1 U544 ( .A1(n533), .A2(n406), .ZN(N2889) );
  NAND2_X1 U545 ( .A1(n442), .A2(n406), .ZN(N2890) );
  INV_X1 U546 ( .A(n406), .ZN(n407) );
  NOR2_X1 U547 ( .A1(n445), .A2(n407), .ZN(N2891) );
  NAND2_X1 U548 ( .A1(n574), .A2(n563), .ZN(n408) );
  NAND2_X1 U549 ( .A1(n556), .A2(n408), .ZN(N2895) );
  NAND2_X1 U550 ( .A1(n446), .A2(n408), .ZN(N2896) );
  INV_X1 U551 ( .A(n408), .ZN(n409) );
  NOR2_X1 U552 ( .A1(n449), .A2(n409), .ZN(N2897) );
  NAND2_X1 U553 ( .A1(n577), .A2(n482), .ZN(n410) );
  NAND2_X1 U554 ( .A1(n471), .A2(n410), .ZN(N2901) );
  NAND2_X1 U555 ( .A1(n434), .A2(n410), .ZN(N2902) );
  INV_X1 U556 ( .A(n410), .ZN(n411) );
  NOR2_X1 U557 ( .A1(n437), .A2(n411), .ZN(N2903) );
  NAND2_X1 U558 ( .A1(n577), .A2(n522), .ZN(n412) );
  NAND2_X1 U559 ( .A1(n517), .A2(n412), .ZN(N2907) );
  NAND2_X1 U560 ( .A1(n438), .A2(n412), .ZN(N2908) );
  INV_X1 U561 ( .A(n412), .ZN(n413) );
  NOR2_X1 U562 ( .A1(n441), .A2(n413), .ZN(N2909) );
  NAND2_X1 U563 ( .A1(n577), .A2(n540), .ZN(n414) );
  NAND2_X1 U564 ( .A1(n533), .A2(n414), .ZN(N2913) );
  NAND2_X1 U565 ( .A1(n442), .A2(n414), .ZN(N2914) );
  INV_X1 U566 ( .A(n414), .ZN(n415) );
  NOR2_X1 U567 ( .A1(n445), .A2(n415), .ZN(N2915) );
  NAND2_X1 U568 ( .A1(n577), .A2(n563), .ZN(n416) );
  NAND2_X1 U569 ( .A1(n556), .A2(n416), .ZN(N2919) );
  NAND2_X1 U570 ( .A1(n446), .A2(n416), .ZN(N2920) );
  INV_X1 U571 ( .A(n416), .ZN(n417) );
  NOR2_X1 U572 ( .A1(n449), .A2(n417), .ZN(N2921) );
  NAND2_X1 U573 ( .A1(n580), .A2(n482), .ZN(n418) );
  NAND2_X1 U574 ( .A1(n471), .A2(n418), .ZN(N2925) );
  NAND2_X1 U575 ( .A1(n434), .A2(n418), .ZN(N2926) );
  INV_X1 U576 ( .A(n418), .ZN(n419) );
  NOR2_X1 U577 ( .A1(n437), .A2(n419), .ZN(N2927) );
  NAND2_X1 U578 ( .A1(n580), .A2(n522), .ZN(n420) );
  NAND2_X1 U579 ( .A1(n517), .A2(n420), .ZN(N2931) );
  NAND2_X1 U580 ( .A1(n438), .A2(n420), .ZN(N2932) );
  INV_X1 U581 ( .A(n420), .ZN(n421) );
  NOR2_X1 U582 ( .A1(n441), .A2(n421), .ZN(N2933) );
  NAND2_X1 U583 ( .A1(n580), .A2(n540), .ZN(n422) );
  NAND2_X1 U584 ( .A1(n533), .A2(n422), .ZN(N2937) );
  NAND2_X1 U585 ( .A1(n442), .A2(n422), .ZN(N2938) );
  INV_X1 U586 ( .A(n422), .ZN(n423) );
  NOR2_X1 U587 ( .A1(n445), .A2(n423), .ZN(N2939) );
  NAND2_X1 U588 ( .A1(n580), .A2(n563), .ZN(n424) );
  NAND2_X1 U589 ( .A1(n556), .A2(n424), .ZN(N2943) );
  NAND2_X1 U590 ( .A1(n446), .A2(n424), .ZN(N2944) );
  INV_X1 U591 ( .A(n424), .ZN(n425) );
  NOR2_X1 U592 ( .A1(n449), .A2(n425), .ZN(N2945) );
  NAND2_X1 U593 ( .A1(n583), .A2(n482), .ZN(n426) );
  NAND2_X1 U594 ( .A1(n471), .A2(n426), .ZN(N2949) );
  NAND2_X1 U595 ( .A1(n434), .A2(n426), .ZN(N2950) );
  INV_X1 U596 ( .A(n426), .ZN(n427) );
  NOR2_X1 U597 ( .A1(n437), .A2(n427), .ZN(N2951) );
  NAND2_X1 U598 ( .A1(n583), .A2(n522), .ZN(n428) );
  NAND2_X1 U599 ( .A1(n517), .A2(n428), .ZN(N2955) );
  NAND2_X1 U600 ( .A1(n438), .A2(n428), .ZN(N2956) );
  INV_X1 U601 ( .A(n428), .ZN(n429) );
  NOR2_X1 U602 ( .A1(n441), .A2(n429), .ZN(N2957) );
  NAND2_X1 U603 ( .A1(n583), .A2(n540), .ZN(n430) );
  NAND2_X1 U604 ( .A1(n533), .A2(n430), .ZN(N2961) );
  NAND2_X1 U605 ( .A1(n442), .A2(n430), .ZN(N2962) );
  INV_X1 U606 ( .A(n430), .ZN(n431) );
  NOR2_X1 U607 ( .A1(n445), .A2(n431), .ZN(N2963) );
  NAND2_X1 U608 ( .A1(n583), .A2(n563), .ZN(n432) );
  NAND2_X1 U609 ( .A1(n556), .A2(n432), .ZN(N2967) );
  NAND2_X1 U610 ( .A1(n446), .A2(n432), .ZN(N2968) );
  INV_X1 U611 ( .A(n432), .ZN(n433) );
  NOR2_X1 U612 ( .A1(n449), .A2(n433), .ZN(N2969) );
  NAND2_X1 U613 ( .A1(n588), .A2(n482), .ZN(n435) );
  NAND2_X1 U614 ( .A1(n471), .A2(n435), .ZN(N2973) );
  NAND2_X1 U615 ( .A1(n434), .A2(n435), .ZN(N2974) );
  INV_X1 U616 ( .A(n435), .ZN(n436) );
  NOR2_X1 U617 ( .A1(n437), .A2(n436), .ZN(N2975) );
  NAND2_X1 U618 ( .A1(n588), .A2(n522), .ZN(n439) );
  NAND2_X1 U619 ( .A1(n517), .A2(n439), .ZN(N2979) );
  NAND2_X1 U620 ( .A1(n438), .A2(n439), .ZN(N2980) );
  INV_X1 U621 ( .A(n439), .ZN(n440) );
  NOR2_X1 U622 ( .A1(n441), .A2(n440), .ZN(N2981) );
  NAND2_X1 U623 ( .A1(n588), .A2(n540), .ZN(n443) );
  NAND2_X1 U624 ( .A1(n533), .A2(n443), .ZN(N2985) );
  NAND2_X1 U625 ( .A1(n442), .A2(n443), .ZN(N2986) );
  INV_X1 U626 ( .A(n443), .ZN(n444) );
  NOR2_X1 U627 ( .A1(n445), .A2(n444), .ZN(N2987) );
  NAND2_X1 U628 ( .A1(n588), .A2(n563), .ZN(n447) );
  NAND2_X1 U629 ( .A1(n556), .A2(n447), .ZN(N2991) );
  NAND2_X1 U630 ( .A1(n446), .A2(n447), .ZN(N2992) );
  INV_X1 U631 ( .A(n447), .ZN(n448) );
  NOR2_X1 U632 ( .A1(n449), .A2(n448), .ZN(N2993) );
  AOI22_X1 U633 ( .A1(n458), .A2(n518), .B1(n455), .B2(n510), .ZN(n450) );
  OAI21_X1 U634 ( .B1(n526), .B2(n460), .A(n450), .ZN(n451) );
  AOI21_X1 U635 ( .B1(n462), .B2(n558), .A(n451), .ZN(n549) );
  AOI22_X1 U636 ( .A1(n458), .A2(n517), .B1(n471), .B2(n510), .ZN(n454) );
  INV_X1 U637 ( .A(n460), .ZN(n452) );
  AOI22_X1 U638 ( .A1(n452), .A2(n533), .B1(n462), .B2(n556), .ZN(n453) );
  NAND2_X1 U639 ( .A1(n454), .A2(n453), .ZN(n546) );
  NOR2_X1 U640 ( .A1(n467), .A2(n546), .ZN(n456) );
  OR2_X1 U641 ( .A1(n456), .A2(n455), .ZN(n457) );
  AOI221_X1 U642 ( .B1(n549), .B2(n457), .C1(n456), .C2(n455), .A(n561), .ZN(
        n466) );
  AOI22_X1 U643 ( .A1(n458), .A2(n514), .B1(n465), .B2(n510), .ZN(n459) );
  OAI21_X1 U644 ( .B1(n536), .B2(n460), .A(n459), .ZN(n461) );
  AOI21_X1 U645 ( .B1(n462), .B2(n553), .A(n461), .ZN(n547) );
  INV_X1 U646 ( .A(n547), .ZN(n535) );
  AOI22_X1 U647 ( .A1(n523), .A2(n514), .B1(n543), .B2(n531), .ZN(n464) );
  NAND2_X1 U648 ( .A1(n564), .A2(n553), .ZN(n463) );
  OAI211_X1 U649 ( .C1(n481), .C2(n474), .A(n464), .B(n463), .ZN(n554) );
  AOI22_X1 U650 ( .A1(n538), .A2(n535), .B1(n554), .B2(n561), .ZN(n552) );
  AOI222_X1 U651 ( .A1(n466), .A2(n465), .B1(n466), .B2(n547), .C1(n465), .C2(
        n552), .ZN(n484) );
  NOR2_X1 U652 ( .A1(n467), .A2(n474), .ZN(n470) );
  AOI221_X1 U653 ( .B1(\last_hit_index[0] ), .B2(n528), .C1(n109), .C2(n468), 
        .A(\last_hit_index[1] ), .ZN(n469) );
  AOI211_X1 U654 ( .C1(n523), .C2(n517), .A(n470), .B(n469), .ZN(n557) );
  NAND2_X1 U655 ( .A1(n557), .A2(n471), .ZN(n476) );
  AOI22_X1 U656 ( .A1(n543), .A2(n534), .B1(n523), .B2(n518), .ZN(n473) );
  NAND2_X1 U657 ( .A1(n564), .A2(n558), .ZN(n472) );
  OAI211_X1 U658 ( .C1(n477), .C2(n474), .A(n473), .B(n472), .ZN(n525) );
  AND2_X1 U659 ( .A1(n477), .A2(n476), .ZN(n475) );
  OAI221_X1 U660 ( .B1(n477), .B2(n476), .C1(n525), .C2(n475), .A(n561), .ZN(
        n478) );
  AOI21_X1 U661 ( .B1(n554), .B2(n481), .A(n478), .ZN(n479) );
  AOI21_X1 U662 ( .B1(n481), .B2(n480), .A(n479), .ZN(n483) );
  NAND2_X1 U663 ( .A1(n509), .A2(n587), .ZN(n565) );
  NOR2_X1 U664 ( .A1(n589), .A2(n565), .ZN(N3093) );
  OAI221_X1 U665 ( .B1(n287), .B2(last_prediction[24]), .C1(n289), .C2(
        last_prediction[25]), .A(n489), .ZN(n496) );
  OAI221_X1 U666 ( .B1(n291), .B2(last_prediction[26]), .C1(n293), .C2(
        last_prediction[27]), .A(n490), .ZN(n495) );
  OAI221_X1 U667 ( .B1(n295), .B2(last_prediction[28]), .C1(n297), .C2(
        last_prediction[29]), .A(n491), .ZN(n494) );
  OAI221_X1 U668 ( .B1(n299), .B2(last_prediction[30]), .C1(n301), .C2(
        last_prediction[31]), .A(n492), .ZN(n493) );
  OAI221_X1 U669 ( .B1(n271), .B2(last_prediction[10]), .C1(n272), .C2(
        last_prediction[11]), .A(n497), .ZN(n503) );
  OAI221_X1 U670 ( .B1(n261), .B2(last_prediction[4]), .C1(n263), .C2(
        last_prediction[5]), .A(n498), .ZN(n501) );
  OAI221_X1 U671 ( .B1(n265), .B2(last_prediction[6]), .C1(n267), .C2(
        last_prediction[7]), .A(n499), .ZN(n500) );
  NOR2_X1 U672 ( .A1(n97), .A2(n565), .ZN(N3094) );
  INV_X1 U673 ( .A(n509), .ZN(n567) );
  NAND3_X1 U674 ( .A1(n538), .A2(n587), .A3(n510), .ZN(n591) );
  NOR2_X1 U675 ( .A1(n567), .A2(n591), .ZN(N3095) );
  OAI21_X1 U676 ( .B1(n549), .B2(n518), .A(n517), .ZN(n511) );
  OAI22_X1 U677 ( .A1(n547), .A2(n514), .B1(n546), .B2(n511), .ZN(n512) );
  AOI211_X1 U678 ( .C1(n549), .C2(n518), .A(n561), .B(n512), .ZN(n513) );
  INV_X1 U679 ( .A(n518), .ZN(n521) );
  AOI21_X1 U680 ( .B1(n516), .B2(n554), .A(n538), .ZN(n520) );
  INV_X1 U681 ( .A(n525), .ZN(n559) );
  OAI211_X1 U682 ( .C1(n559), .C2(n518), .A(n557), .B(n517), .ZN(n519) );
  NOR2_X1 U683 ( .A1(n592), .A2(n565), .ZN(N3096) );
  NOR2_X1 U684 ( .A1(n565), .A2(n102), .ZN(N3097) );
  NOR2_X1 U685 ( .A1(n567), .A2(n594), .ZN(N3098) );
  OAI21_X1 U686 ( .B1(n559), .B2(n534), .A(n557), .ZN(n527) );
  OAI22_X1 U687 ( .A1(n528), .A2(n527), .B1(n526), .B2(n525), .ZN(n529) );
  AOI211_X1 U688 ( .C1(n536), .C2(n554), .A(n538), .B(n529), .ZN(n530) );
  AOI221_X1 U689 ( .B1(n532), .B2(n536), .C1(n552), .C2(n531), .A(n530), .ZN(
        n542) );
  OAI21_X1 U690 ( .B1(n549), .B2(n534), .A(n533), .ZN(n539) );
  AOI22_X1 U691 ( .A1(n536), .A2(n535), .B1(n549), .B2(n534), .ZN(n537) );
  OAI211_X1 U692 ( .C1(n539), .C2(n546), .A(n538), .B(n537), .ZN(n541) );
  NOR2_X1 U693 ( .A1(n595), .A2(n565), .ZN(N3099) );
  NOR2_X1 U694 ( .A1(n565), .A2(n103), .ZN(N3100) );
  NOR2_X1 U695 ( .A1(n567), .A2(n597), .ZN(N3101) );
  OAI21_X1 U696 ( .B1(n549), .B2(n558), .A(n556), .ZN(n545) );
  OAI22_X1 U697 ( .A1(n547), .A2(n553), .B1(n546), .B2(n545), .ZN(n548) );
  AOI211_X1 U698 ( .C1(n549), .C2(n558), .A(n561), .B(n548), .ZN(n551) );
  AOI22_X1 U699 ( .A1(n555), .A2(n554), .B1(n559), .B2(n558), .ZN(n562) );
  OAI211_X1 U700 ( .C1(n559), .C2(n558), .A(n557), .B(n556), .ZN(n560) );
  NOR2_X1 U701 ( .A1(n598), .A2(n565), .ZN(N3102) );
  NOR2_X1 U702 ( .A1(n565), .A2(n99), .ZN(N3103) );
  NOR2_X1 U703 ( .A1(n567), .A2(n601), .ZN(N3104) );
  NAND2_X1 U704 ( .A1(n568), .A2(n587), .ZN(n569) );
  NOR2_X1 U705 ( .A1(n589), .A2(n569), .ZN(N3105) );
  NOR2_X1 U706 ( .A1(n97), .A2(n569), .ZN(N3106) );
  NOR2_X1 U707 ( .A1(n570), .A2(n591), .ZN(N3107) );
  NOR2_X1 U708 ( .A1(n592), .A2(n569), .ZN(N3108) );
  NOR2_X1 U709 ( .A1(n101), .A2(n569), .ZN(N3109) );
  NOR2_X1 U710 ( .A1(n570), .A2(n594), .ZN(N3110) );
  NOR2_X1 U711 ( .A1(n595), .A2(n569), .ZN(N3111) );
  NOR2_X1 U712 ( .A1(n569), .A2(n103), .ZN(N3112) );
  NOR2_X1 U713 ( .A1(n570), .A2(n597), .ZN(N3113) );
  NOR2_X1 U714 ( .A1(n598), .A2(n569), .ZN(N3114) );
  NOR2_X1 U715 ( .A1(n569), .A2(n99), .ZN(N3115) );
  NOR2_X1 U716 ( .A1(n570), .A2(n601), .ZN(N3116) );
  NAND2_X1 U717 ( .A1(n571), .A2(n587), .ZN(n572) );
  NOR2_X1 U718 ( .A1(n589), .A2(n572), .ZN(N3117) );
  NOR2_X1 U719 ( .A1(n97), .A2(n572), .ZN(N3118) );
  INV_X1 U720 ( .A(n571), .ZN(n573) );
  NOR2_X1 U721 ( .A1(n573), .A2(n591), .ZN(N3119) );
  NOR2_X1 U722 ( .A1(n592), .A2(n572), .ZN(N3120) );
  NOR2_X1 U723 ( .A1(n572), .A2(n102), .ZN(N3121) );
  NOR2_X1 U724 ( .A1(n573), .A2(n594), .ZN(N3122) );
  NOR2_X1 U725 ( .A1(n595), .A2(n572), .ZN(N3123) );
  NOR2_X1 U726 ( .A1(n572), .A2(n103), .ZN(N3124) );
  NOR2_X1 U727 ( .A1(n573), .A2(n597), .ZN(N3125) );
  NOR2_X1 U728 ( .A1(n598), .A2(n572), .ZN(N3126) );
  NOR2_X1 U729 ( .A1(n572), .A2(n99), .ZN(N3127) );
  NOR2_X1 U730 ( .A1(n573), .A2(n601), .ZN(N3128) );
  NAND2_X1 U731 ( .A1(n574), .A2(n587), .ZN(n575) );
  NOR2_X1 U732 ( .A1(n589), .A2(n575), .ZN(N3129) );
  NOR2_X1 U733 ( .A1(n98), .A2(n575), .ZN(N3130) );
  NOR2_X1 U734 ( .A1(n576), .A2(n591), .ZN(N3131) );
  NOR2_X1 U735 ( .A1(n592), .A2(n575), .ZN(N3132) );
  NOR2_X1 U736 ( .A1(n575), .A2(n101), .ZN(N3133) );
  NOR2_X1 U737 ( .A1(n576), .A2(n594), .ZN(N3134) );
  NOR2_X1 U738 ( .A1(n595), .A2(n575), .ZN(N3135) );
  NOR2_X1 U739 ( .A1(n575), .A2(n104), .ZN(N3136) );
  NOR2_X1 U740 ( .A1(n576), .A2(n597), .ZN(N3137) );
  NOR2_X1 U741 ( .A1(n598), .A2(n575), .ZN(N3138) );
  NOR2_X1 U742 ( .A1(n575), .A2(n100), .ZN(N3139) );
  NOR2_X1 U743 ( .A1(n576), .A2(n601), .ZN(N3140) );
  NAND2_X1 U744 ( .A1(n577), .A2(n587), .ZN(n578) );
  NOR2_X1 U745 ( .A1(n589), .A2(n578), .ZN(N3141) );
  NOR2_X1 U746 ( .A1(n98), .A2(n578), .ZN(N3142) );
  NOR2_X1 U747 ( .A1(n579), .A2(n591), .ZN(N3143) );
  NOR2_X1 U748 ( .A1(n592), .A2(n578), .ZN(N3144) );
  NOR2_X1 U749 ( .A1(n578), .A2(n102), .ZN(N3145) );
  NOR2_X1 U750 ( .A1(n579), .A2(n594), .ZN(N3146) );
  NOR2_X1 U751 ( .A1(n595), .A2(n578), .ZN(N3147) );
  NOR2_X1 U752 ( .A1(n578), .A2(n104), .ZN(N3148) );
  NOR2_X1 U753 ( .A1(n579), .A2(n597), .ZN(N3149) );
  NOR2_X1 U754 ( .A1(n598), .A2(n578), .ZN(N3150) );
  NOR2_X1 U755 ( .A1(n578), .A2(n100), .ZN(N3151) );
  NOR2_X1 U756 ( .A1(n579), .A2(n601), .ZN(N3152) );
  NAND2_X1 U757 ( .A1(n580), .A2(n587), .ZN(n581) );
  NOR2_X1 U758 ( .A1(n589), .A2(n581), .ZN(N3153) );
  NOR2_X1 U759 ( .A1(n98), .A2(n581), .ZN(N3154) );
  NOR2_X1 U760 ( .A1(n582), .A2(n591), .ZN(N3155) );
  NOR2_X1 U761 ( .A1(n592), .A2(n581), .ZN(N3156) );
  NOR2_X1 U762 ( .A1(n581), .A2(n101), .ZN(N3157) );
  NOR2_X1 U763 ( .A1(n582), .A2(n594), .ZN(N3158) );
  NOR2_X1 U764 ( .A1(n595), .A2(n581), .ZN(N3159) );
  NOR2_X1 U765 ( .A1(n581), .A2(n104), .ZN(N3160) );
  NOR2_X1 U766 ( .A1(n582), .A2(n597), .ZN(N3161) );
  NOR2_X1 U767 ( .A1(n598), .A2(n581), .ZN(N3162) );
  NOR2_X1 U768 ( .A1(n581), .A2(n100), .ZN(N3163) );
  NOR2_X1 U769 ( .A1(n582), .A2(n601), .ZN(N3164) );
  NAND2_X1 U770 ( .A1(n583), .A2(n587), .ZN(n584) );
  NOR2_X1 U771 ( .A1(n589), .A2(n584), .ZN(N3165) );
  NOR2_X1 U772 ( .A1(n97), .A2(n584), .ZN(N3166) );
  NOR2_X1 U773 ( .A1(n586), .A2(n591), .ZN(N3167) );
  NOR2_X1 U774 ( .A1(n592), .A2(n584), .ZN(N3168) );
  NOR2_X1 U775 ( .A1(n584), .A2(n102), .ZN(N3169) );
  NOR2_X1 U776 ( .A1(n586), .A2(n594), .ZN(N3170) );
  NOR2_X1 U777 ( .A1(n595), .A2(n584), .ZN(N3171) );
  NOR2_X1 U778 ( .A1(n584), .A2(n103), .ZN(N3172) );
  NOR2_X1 U779 ( .A1(n586), .A2(n597), .ZN(N3173) );
  NOR2_X1 U780 ( .A1(n598), .A2(n584), .ZN(N3174) );
  NOR2_X1 U781 ( .A1(n584), .A2(n99), .ZN(N3175) );
  NOR2_X1 U782 ( .A1(n586), .A2(n601), .ZN(N3176) );
  NAND2_X1 U783 ( .A1(n588), .A2(n587), .ZN(n600) );
  NOR2_X1 U784 ( .A1(n589), .A2(n600), .ZN(N3177) );
  NOR2_X1 U785 ( .A1(n98), .A2(n600), .ZN(N3178) );
  NOR2_X1 U786 ( .A1(n602), .A2(n591), .ZN(N3179) );
  NOR2_X1 U787 ( .A1(n592), .A2(n600), .ZN(N3180) );
  NOR2_X1 U788 ( .A1(n600), .A2(n101), .ZN(N3181) );
  NOR2_X1 U789 ( .A1(n602), .A2(n594), .ZN(N3182) );
  NOR2_X1 U790 ( .A1(n595), .A2(n600), .ZN(N3183) );
  NOR2_X1 U791 ( .A1(n600), .A2(n104), .ZN(N3184) );
  NOR2_X1 U792 ( .A1(n602), .A2(n597), .ZN(N3185) );
  NOR2_X1 U793 ( .A1(n598), .A2(n600), .ZN(N3186) );
  NOR2_X1 U794 ( .A1(n600), .A2(n100), .ZN(N3187) );
  NOR2_X1 U795 ( .A1(n602), .A2(n601), .ZN(N3188) );
  INV_X1 U796 ( .A(instr_fetch[28]), .ZN(n604) );
  NOR3_X1 U797 ( .A1(instr_fetch[27]), .A2(n604), .A3(instr_fetch[30]), .ZN(
        n603) );
  AOI21_X1 U798 ( .B1(n604), .B2(instr_fetch[27]), .A(n603), .ZN(n605) );
  NOR3_X1 U799 ( .A1(instr_fetch[29]), .A2(instr_fetch[31]), .A3(n605), .ZN(
        n906) );
  NAND2_X1 U800 ( .A1(n882), .A2(IF_EN), .ZN(n606) );
  INV_X1 U801 ( .A(n606), .ZN(N3361) );
  INV_X1 U802 ( .A(pc_fetch[6]), .ZN(n67) );
  INV_X1 U803 ( .A(pc_fetch[12]), .ZN(n64) );
  NOR3_X1 U804 ( .A1(pc_fetch[2]), .A2(n1586), .A3(n608), .ZN(n1569) );
  NOR3_X1 U805 ( .A1(n609), .A2(n1586), .A3(n608), .ZN(n1568) );
  AOI22_X1 U806 ( .A1(n57), .A2(\cache[0][0][TAG][4] ), .B1(n36), .B2(
        \cache[1][0][TAG][4] ), .ZN(n613) );
  AOI22_X1 U807 ( .A1(n240), .A2(\cache[2][0][TAG][4] ), .B1(n37), .B2(
        \cache[3][0][TAG][4] ), .ZN(n612) );
  AOI22_X1 U808 ( .A1(n244), .A2(\cache[4][0][TAG][4] ), .B1(n38), .B2(
        \cache[5][0][TAG][4] ), .ZN(n611) );
  NOR3_X1 U809 ( .A1(pc_fetch[2]), .A2(pc_fetch[3]), .A3(pc_fetch[4]), .ZN(
        n1575) );
  NOR3_X1 U810 ( .A1(pc_fetch[3]), .A2(pc_fetch[4]), .A3(n609), .ZN(n1574) );
  AOI22_X1 U811 ( .A1(n40), .A2(\cache[6][0][TAG][4] ), .B1(n39), .B2(
        \cache[7][0][TAG][4] ), .ZN(n610) );
  AND4_X1 U812 ( .A1(n613), .A2(n612), .A3(n611), .A4(n610), .ZN(n620) );
  INV_X1 U813 ( .A(pc_fetch[11]), .ZN(n750) );
  AOI22_X1 U814 ( .A1(n57), .A2(\cache[0][0][TAG][6] ), .B1(n232), .B2(
        \cache[1][0][TAG][6] ), .ZN(n617) );
  AOI22_X1 U815 ( .A1(n55), .A2(\cache[2][0][TAG][6] ), .B1(n238), .B2(
        \cache[3][0][TAG][6] ), .ZN(n616) );
  AOI22_X1 U816 ( .A1(n56), .A2(\cache[4][0][TAG][6] ), .B1(n242), .B2(
        \cache[5][0][TAG][6] ), .ZN(n615) );
  AOI22_X1 U817 ( .A1(n40), .A2(\cache[6][0][TAG][6] ), .B1(n246), .B2(
        \cache[7][0][TAG][6] ), .ZN(n614) );
  NAND4_X1 U818 ( .A1(n617), .A2(n616), .A3(n615), .A4(n614), .ZN(n619) );
  AOI22_X1 U819 ( .A1(pc_fetch[9]), .A2(n620), .B1(n619), .B2(n750), .ZN(n618)
         );
  OAI221_X1 U820 ( .B1(pc_fetch[9]), .B2(n620), .C1(n750), .C2(n619), .A(n618), 
        .ZN(n674) );
  AOI22_X1 U821 ( .A1(n57), .A2(\cache[0][0][TAG][7] ), .B1(n232), .B2(
        \cache[1][0][TAG][7] ), .ZN(n624) );
  AOI22_X1 U822 ( .A1(n239), .A2(\cache[2][0][TAG][7] ), .B1(n238), .B2(
        \cache[3][0][TAG][7] ), .ZN(n623) );
  AOI22_X1 U823 ( .A1(n243), .A2(\cache[4][0][TAG][7] ), .B1(n242), .B2(
        \cache[5][0][TAG][7] ), .ZN(n622) );
  AOI22_X1 U824 ( .A1(n40), .A2(\cache[6][0][TAG][7] ), .B1(n246), .B2(
        \cache[7][0][TAG][7] ), .ZN(n621) );
  AND4_X1 U825 ( .A1(n624), .A2(n623), .A3(n622), .A4(n621), .ZN(n631) );
  AOI22_X1 U826 ( .A1(n57), .A2(\cache[0][0][TAG][5] ), .B1(n232), .B2(
        \cache[1][0][TAG][5] ), .ZN(n628) );
  AOI22_X1 U827 ( .A1(n239), .A2(\cache[2][0][TAG][5] ), .B1(n238), .B2(
        \cache[3][0][TAG][5] ), .ZN(n627) );
  AOI22_X1 U828 ( .A1(n243), .A2(\cache[4][0][TAG][5] ), .B1(n242), .B2(
        \cache[5][0][TAG][5] ), .ZN(n626) );
  AOI22_X1 U829 ( .A1(n40), .A2(\cache[6][0][TAG][5] ), .B1(n246), .B2(
        \cache[7][0][TAG][5] ), .ZN(n625) );
  NAND4_X1 U830 ( .A1(n628), .A2(n627), .A3(n626), .A4(n625), .ZN(n630) );
  AOI22_X1 U831 ( .A1(pc_fetch[12]), .A2(n631), .B1(n630), .B2(n65), .ZN(n629)
         );
  OAI221_X1 U832 ( .B1(pc_fetch[12]), .B2(n631), .C1(n65), .C2(n630), .A(n629), 
        .ZN(n673) );
  AOI22_X1 U833 ( .A1(n57), .A2(\cache[0][0][TAG][1] ), .B1(n232), .B2(
        \cache[1][0][TAG][1] ), .ZN(n635) );
  AOI22_X1 U834 ( .A1(n239), .A2(\cache[2][0][TAG][1] ), .B1(n238), .B2(
        \cache[3][0][TAG][1] ), .ZN(n634) );
  AOI22_X1 U835 ( .A1(n243), .A2(\cache[4][0][TAG][1] ), .B1(n242), .B2(
        \cache[5][0][TAG][1] ), .ZN(n633) );
  AOI22_X1 U836 ( .A1(n40), .A2(\cache[6][0][TAG][1] ), .B1(n246), .B2(
        \cache[7][0][TAG][1] ), .ZN(n632) );
  AND4_X1 U837 ( .A1(n635), .A2(n634), .A3(n633), .A4(n632), .ZN(n642) );
  AOI22_X1 U838 ( .A1(n57), .A2(\cache[0][0][TAG][3] ), .B1(n232), .B2(
        \cache[1][0][TAG][3] ), .ZN(n639) );
  AOI22_X1 U839 ( .A1(n239), .A2(\cache[2][0][TAG][3] ), .B1(n238), .B2(
        \cache[3][0][TAG][3] ), .ZN(n638) );
  AOI22_X1 U840 ( .A1(n243), .A2(\cache[4][0][TAG][3] ), .B1(n242), .B2(
        \cache[5][0][TAG][3] ), .ZN(n637) );
  AOI22_X1 U841 ( .A1(n40), .A2(\cache[6][0][TAG][3] ), .B1(n246), .B2(
        \cache[7][0][TAG][3] ), .ZN(n636) );
  NAND4_X1 U842 ( .A1(n639), .A2(n638), .A3(n637), .A4(n636), .ZN(n641) );
  AOI22_X1 U843 ( .A1(pc_fetch[6]), .A2(n642), .B1(n641), .B2(n66), .ZN(n640)
         );
  OAI221_X1 U844 ( .B1(pc_fetch[6]), .B2(n642), .C1(n66), .C2(n641), .A(n640), 
        .ZN(n672) );
  AOI22_X1 U845 ( .A1(\cache[0][0][YOUTH][2] ), .A2(n57), .B1(
        \cache[1][0][YOUTH][2] ), .B2(n36), .ZN(n646) );
  AOI22_X1 U846 ( .A1(\cache[3][0][YOUTH][2] ), .A2(n37), .B1(
        \cache[2][0][YOUTH][2] ), .B2(n240), .ZN(n645) );
  AOI22_X1 U847 ( .A1(\cache[5][0][YOUTH][2] ), .A2(n38), .B1(
        \cache[4][0][YOUTH][2] ), .B2(n244), .ZN(n644) );
  AOI22_X1 U848 ( .A1(\cache[7][0][YOUTH][2] ), .A2(n39), .B1(
        \cache[6][0][YOUTH][2] ), .B2(n40), .ZN(n643) );
  NAND4_X1 U849 ( .A1(n646), .A2(n645), .A3(n644), .A4(n643), .ZN(n657) );
  AOI22_X1 U850 ( .A1(\cache[0][0][YOUTH][0] ), .A2(n57), .B1(
        \cache[1][0][YOUTH][0] ), .B2(n36), .ZN(n650) );
  AOI22_X1 U851 ( .A1(\cache[3][0][YOUTH][0] ), .A2(n37), .B1(
        \cache[2][0][YOUTH][0] ), .B2(n55), .ZN(n649) );
  AOI22_X1 U852 ( .A1(\cache[5][0][YOUTH][0] ), .A2(n38), .B1(
        \cache[4][0][YOUTH][0] ), .B2(n56), .ZN(n648) );
  AOI22_X1 U853 ( .A1(\cache[7][0][YOUTH][0] ), .A2(n39), .B1(
        \cache[6][0][YOUTH][0] ), .B2(n40), .ZN(n647) );
  NAND4_X1 U854 ( .A1(n650), .A2(n649), .A3(n648), .A4(n647), .ZN(n656) );
  AOI22_X1 U855 ( .A1(\cache[0][0][YOUTH][1] ), .A2(n57), .B1(
        \cache[1][0][YOUTH][1] ), .B2(n36), .ZN(n654) );
  AOI22_X1 U856 ( .A1(\cache[3][0][YOUTH][1] ), .A2(n37), .B1(
        \cache[2][0][YOUTH][1] ), .B2(n239), .ZN(n653) );
  AOI22_X1 U857 ( .A1(\cache[5][0][YOUTH][1] ), .A2(n38), .B1(
        \cache[4][0][YOUTH][1] ), .B2(n243), .ZN(n652) );
  AOI22_X1 U858 ( .A1(\cache[7][0][YOUTH][1] ), .A2(n39), .B1(
        \cache[6][0][YOUTH][1] ), .B2(n40), .ZN(n651) );
  NAND4_X1 U859 ( .A1(n654), .A2(n653), .A3(n652), .A4(n651), .ZN(n655) );
  NAND3_X1 U860 ( .A1(n657), .A2(n656), .A3(n655), .ZN(n670) );
  AOI22_X1 U861 ( .A1(n57), .A2(\cache[0][0][TAG][0] ), .B1(n232), .B2(
        \cache[1][0][TAG][0] ), .ZN(n661) );
  AOI22_X1 U862 ( .A1(n240), .A2(\cache[2][0][TAG][0] ), .B1(n238), .B2(
        \cache[3][0][TAG][0] ), .ZN(n660) );
  AOI22_X1 U863 ( .A1(n244), .A2(\cache[4][0][TAG][0] ), .B1(n242), .B2(
        \cache[5][0][TAG][0] ), .ZN(n659) );
  AOI22_X1 U864 ( .A1(n40), .A2(\cache[6][0][TAG][0] ), .B1(n246), .B2(
        \cache[7][0][TAG][0] ), .ZN(n658) );
  NAND4_X1 U865 ( .A1(n661), .A2(n660), .A3(n659), .A4(n658), .ZN(n668) );
  INV_X1 U866 ( .A(pc_fetch[5]), .ZN(n799) );
  AOI22_X1 U867 ( .A1(n57), .A2(\cache[0][0][TAG][2] ), .B1(n232), .B2(
        \cache[1][0][TAG][2] ), .ZN(n665) );
  AOI22_X1 U868 ( .A1(n240), .A2(\cache[2][0][TAG][2] ), .B1(n238), .B2(
        \cache[3][0][TAG][2] ), .ZN(n664) );
  AOI22_X1 U869 ( .A1(n244), .A2(\cache[4][0][TAG][2] ), .B1(n242), .B2(
        \cache[5][0][TAG][2] ), .ZN(n663) );
  AOI22_X1 U870 ( .A1(n40), .A2(\cache[6][0][TAG][2] ), .B1(n246), .B2(
        \cache[7][0][TAG][2] ), .ZN(n662) );
  AND4_X1 U871 ( .A1(n665), .A2(n664), .A3(n663), .A4(n662), .ZN(n667) );
  OAI22_X1 U872 ( .A1(n799), .A2(n668), .B1(pc_fetch[7]), .B2(n667), .ZN(n666)
         );
  AOI221_X1 U873 ( .B1(n668), .B2(n799), .C1(pc_fetch[7]), .C2(n667), .A(n666), 
        .ZN(n669) );
  NAND2_X1 U874 ( .A1(n670), .A2(n669), .ZN(n671) );
  NOR4_X1 U875 ( .A1(n674), .A2(n673), .A3(n672), .A4(n671), .ZN(n807) );
  AOI22_X1 U876 ( .A1(n57), .A2(\cache[0][1][TAG][0] ), .B1(n232), .B2(
        \cache[1][1][TAG][0] ), .ZN(n678) );
  AOI22_X1 U877 ( .A1(n239), .A2(\cache[2][1][TAG][0] ), .B1(n238), .B2(
        \cache[3][1][TAG][0] ), .ZN(n677) );
  AOI22_X1 U878 ( .A1(n243), .A2(\cache[4][1][TAG][0] ), .B1(n242), .B2(
        \cache[5][1][TAG][0] ), .ZN(n676) );
  AOI22_X1 U879 ( .A1(n40), .A2(\cache[6][1][TAG][0] ), .B1(n246), .B2(
        \cache[7][1][TAG][0] ), .ZN(n675) );
  NAND4_X1 U880 ( .A1(n678), .A2(n677), .A3(n676), .A4(n675), .ZN(n685) );
  AOI22_X1 U881 ( .A1(n57), .A2(\cache[0][1][TAG][2] ), .B1(n232), .B2(
        \cache[1][1][TAG][2] ), .ZN(n682) );
  AOI22_X1 U882 ( .A1(n239), .A2(\cache[2][1][TAG][2] ), .B1(n238), .B2(
        \cache[3][1][TAG][2] ), .ZN(n681) );
  AOI22_X1 U883 ( .A1(n243), .A2(\cache[4][1][TAG][2] ), .B1(n242), .B2(
        \cache[5][1][TAG][2] ), .ZN(n680) );
  AOI22_X1 U884 ( .A1(n40), .A2(\cache[6][1][TAG][2] ), .B1(n246), .B2(
        \cache[7][1][TAG][2] ), .ZN(n679) );
  AND4_X1 U885 ( .A1(n682), .A2(n681), .A3(n680), .A4(n679), .ZN(n684) );
  OAI22_X1 U886 ( .A1(n799), .A2(n685), .B1(pc_fetch[7]), .B2(n684), .ZN(n683)
         );
  AOI221_X1 U887 ( .B1(n685), .B2(n799), .C1(pc_fetch[7]), .C2(n684), .A(n683), 
        .ZN(n739) );
  AOI22_X1 U888 ( .A1(n57), .A2(\cache[0][1][TAG][4] ), .B1(n232), .B2(
        \cache[1][1][TAG][4] ), .ZN(n689) );
  AOI22_X1 U889 ( .A1(n55), .A2(\cache[2][1][TAG][4] ), .B1(n238), .B2(
        \cache[3][1][TAG][4] ), .ZN(n688) );
  AOI22_X1 U890 ( .A1(n56), .A2(\cache[4][1][TAG][4] ), .B1(n242), .B2(
        \cache[5][1][TAG][4] ), .ZN(n687) );
  AOI22_X1 U891 ( .A1(n40), .A2(\cache[6][1][TAG][4] ), .B1(n246), .B2(
        \cache[7][1][TAG][4] ), .ZN(n686) );
  AND4_X1 U892 ( .A1(n689), .A2(n688), .A3(n687), .A4(n686), .ZN(n696) );
  AOI22_X1 U893 ( .A1(n234), .A2(\cache[0][1][TAG][6] ), .B1(n36), .B2(
        \cache[1][1][TAG][6] ), .ZN(n693) );
  AOI22_X1 U894 ( .A1(n239), .A2(\cache[2][1][TAG][6] ), .B1(n37), .B2(
        \cache[3][1][TAG][6] ), .ZN(n692) );
  AOI22_X1 U895 ( .A1(n243), .A2(\cache[4][1][TAG][6] ), .B1(n38), .B2(
        \cache[5][1][TAG][6] ), .ZN(n691) );
  AOI22_X1 U896 ( .A1(n40), .A2(\cache[6][1][TAG][6] ), .B1(n39), .B2(
        \cache[7][1][TAG][6] ), .ZN(n690) );
  NAND4_X1 U897 ( .A1(n693), .A2(n692), .A3(n691), .A4(n690), .ZN(n695) );
  AOI22_X1 U898 ( .A1(pc_fetch[9]), .A2(n696), .B1(n695), .B2(n750), .ZN(n694)
         );
  OAI221_X1 U899 ( .B1(pc_fetch[9]), .B2(n696), .C1(n750), .C2(n695), .A(n694), 
        .ZN(n721) );
  AOI22_X1 U900 ( .A1(n57), .A2(\cache[0][1][TAG][7] ), .B1(n36), .B2(
        \cache[1][1][TAG][7] ), .ZN(n700) );
  AOI22_X1 U901 ( .A1(n55), .A2(\cache[2][1][TAG][7] ), .B1(n37), .B2(
        \cache[3][1][TAG][7] ), .ZN(n699) );
  AOI22_X1 U902 ( .A1(n56), .A2(\cache[4][1][TAG][7] ), .B1(n38), .B2(
        \cache[5][1][TAG][7] ), .ZN(n698) );
  AOI22_X1 U903 ( .A1(n40), .A2(\cache[6][1][TAG][7] ), .B1(n39), .B2(
        \cache[7][1][TAG][7] ), .ZN(n697) );
  AND4_X1 U904 ( .A1(n700), .A2(n699), .A3(n698), .A4(n697), .ZN(n707) );
  AOI22_X1 U905 ( .A1(n234), .A2(\cache[0][1][TAG][5] ), .B1(n36), .B2(
        \cache[1][1][TAG][5] ), .ZN(n704) );
  AOI22_X1 U906 ( .A1(n55), .A2(\cache[2][1][TAG][5] ), .B1(n37), .B2(
        \cache[3][1][TAG][5] ), .ZN(n703) );
  AOI22_X1 U907 ( .A1(n56), .A2(\cache[4][1][TAG][5] ), .B1(n38), .B2(
        \cache[5][1][TAG][5] ), .ZN(n702) );
  AOI22_X1 U908 ( .A1(n40), .A2(\cache[6][1][TAG][5] ), .B1(n39), .B2(
        \cache[7][1][TAG][5] ), .ZN(n701) );
  NAND4_X1 U909 ( .A1(n704), .A2(n703), .A3(n702), .A4(n701), .ZN(n706) );
  AOI22_X1 U910 ( .A1(pc_fetch[12]), .A2(n707), .B1(n706), .B2(n65), .ZN(n705)
         );
  OAI221_X1 U911 ( .B1(pc_fetch[12]), .B2(n707), .C1(n65), .C2(n706), .A(n705), 
        .ZN(n720) );
  AOI22_X1 U912 ( .A1(n57), .A2(\cache[0][1][TAG][1] ), .B1(n36), .B2(
        \cache[1][1][TAG][1] ), .ZN(n711) );
  AOI22_X1 U913 ( .A1(n55), .A2(\cache[2][1][TAG][1] ), .B1(n37), .B2(
        \cache[3][1][TAG][1] ), .ZN(n710) );
  AOI22_X1 U914 ( .A1(n56), .A2(\cache[4][1][TAG][1] ), .B1(n38), .B2(
        \cache[5][1][TAG][1] ), .ZN(n709) );
  AOI22_X1 U915 ( .A1(n40), .A2(\cache[6][1][TAG][1] ), .B1(n39), .B2(
        \cache[7][1][TAG][1] ), .ZN(n708) );
  AND4_X1 U916 ( .A1(n711), .A2(n710), .A3(n709), .A4(n708), .ZN(n718) );
  AOI22_X1 U917 ( .A1(n234), .A2(\cache[0][1][TAG][3] ), .B1(n36), .B2(
        \cache[1][1][TAG][3] ), .ZN(n715) );
  AOI22_X1 U918 ( .A1(n55), .A2(\cache[2][1][TAG][3] ), .B1(n37), .B2(
        \cache[3][1][TAG][3] ), .ZN(n714) );
  AOI22_X1 U919 ( .A1(n56), .A2(\cache[4][1][TAG][3] ), .B1(n38), .B2(
        \cache[5][1][TAG][3] ), .ZN(n713) );
  AOI22_X1 U920 ( .A1(n40), .A2(\cache[6][1][TAG][3] ), .B1(n39), .B2(
        \cache[7][1][TAG][3] ), .ZN(n712) );
  NAND4_X1 U921 ( .A1(n715), .A2(n714), .A3(n713), .A4(n712), .ZN(n717) );
  AOI22_X1 U922 ( .A1(pc_fetch[6]), .A2(n718), .B1(n717), .B2(n66), .ZN(n716)
         );
  OAI221_X1 U923 ( .B1(pc_fetch[6]), .B2(n718), .C1(n66), .C2(n717), .A(n716), 
        .ZN(n719) );
  NOR3_X1 U924 ( .A1(n721), .A2(n720), .A3(n719), .ZN(n738) );
  AOI22_X1 U925 ( .A1(\cache[0][1][YOUTH][1] ), .A2(n57), .B1(
        \cache[1][1][YOUTH][1] ), .B2(n36), .ZN(n725) );
  AOI22_X1 U926 ( .A1(\cache[3][1][YOUTH][1] ), .A2(n37), .B1(
        \cache[2][1][YOUTH][1] ), .B2(n240), .ZN(n724) );
  AOI22_X1 U927 ( .A1(\cache[5][1][YOUTH][1] ), .A2(n38), .B1(
        \cache[4][1][YOUTH][1] ), .B2(n244), .ZN(n723) );
  AOI22_X1 U928 ( .A1(\cache[7][1][YOUTH][1] ), .A2(n39), .B1(
        \cache[6][1][YOUTH][1] ), .B2(n40), .ZN(n722) );
  NAND4_X1 U929 ( .A1(n725), .A2(n724), .A3(n723), .A4(n722), .ZN(n736) );
  AOI22_X1 U930 ( .A1(\cache[0][1][YOUTH][2] ), .A2(n57), .B1(
        \cache[1][1][YOUTH][2] ), .B2(n36), .ZN(n729) );
  AOI22_X1 U931 ( .A1(\cache[3][1][YOUTH][2] ), .A2(n37), .B1(
        \cache[2][1][YOUTH][2] ), .B2(n1571), .ZN(n728) );
  AOI22_X1 U932 ( .A1(\cache[5][1][YOUTH][2] ), .A2(n38), .B1(
        \cache[4][1][YOUTH][2] ), .B2(n1573), .ZN(n727) );
  AOI22_X1 U933 ( .A1(\cache[7][1][YOUTH][2] ), .A2(n39), .B1(
        \cache[6][1][YOUTH][2] ), .B2(n40), .ZN(n726) );
  NAND4_X1 U934 ( .A1(n729), .A2(n728), .A3(n727), .A4(n726), .ZN(n735) );
  AOI22_X1 U935 ( .A1(\cache[0][1][YOUTH][0] ), .A2(n57), .B1(
        \cache[1][1][YOUTH][0] ), .B2(n36), .ZN(n733) );
  AOI22_X1 U936 ( .A1(\cache[3][1][YOUTH][0] ), .A2(n37), .B1(
        \cache[2][1][YOUTH][0] ), .B2(n1571), .ZN(n732) );
  AOI22_X1 U937 ( .A1(\cache[5][1][YOUTH][0] ), .A2(n38), .B1(
        \cache[4][1][YOUTH][0] ), .B2(n1573), .ZN(n731) );
  AOI22_X1 U938 ( .A1(\cache[7][1][YOUTH][0] ), .A2(n39), .B1(
        \cache[6][1][YOUTH][0] ), .B2(n40), .ZN(n730) );
  NAND4_X1 U939 ( .A1(n733), .A2(n732), .A3(n731), .A4(n730), .ZN(n734) );
  NAND3_X1 U940 ( .A1(n736), .A2(n735), .A3(n734), .ZN(n737) );
  NAND3_X1 U941 ( .A1(n739), .A2(n738), .A3(n737), .ZN(n884) );
  AOI22_X1 U942 ( .A1(n234), .A2(\cache[0][2][TAG][4] ), .B1(n36), .B2(
        \cache[1][2][TAG][4] ), .ZN(n743) );
  AOI22_X1 U943 ( .A1(n55), .A2(\cache[2][2][TAG][4] ), .B1(n37), .B2(
        \cache[3][2][TAG][4] ), .ZN(n742) );
  AOI22_X1 U944 ( .A1(n56), .A2(\cache[4][2][TAG][4] ), .B1(n38), .B2(
        \cache[5][2][TAG][4] ), .ZN(n741) );
  AOI22_X1 U945 ( .A1(n40), .A2(\cache[6][2][TAG][4] ), .B1(n39), .B2(
        \cache[7][2][TAG][4] ), .ZN(n740) );
  AND4_X1 U946 ( .A1(n743), .A2(n742), .A3(n741), .A4(n740), .ZN(n751) );
  AOI22_X1 U947 ( .A1(n236), .A2(\cache[0][2][TAG][6] ), .B1(n36), .B2(
        \cache[1][2][TAG][6] ), .ZN(n747) );
  AOI22_X1 U948 ( .A1(n239), .A2(\cache[2][2][TAG][6] ), .B1(n37), .B2(
        \cache[3][2][TAG][6] ), .ZN(n746) );
  AOI22_X1 U949 ( .A1(n243), .A2(\cache[4][2][TAG][6] ), .B1(n38), .B2(
        \cache[5][2][TAG][6] ), .ZN(n745) );
  AOI22_X1 U950 ( .A1(n40), .A2(\cache[6][2][TAG][6] ), .B1(n39), .B2(
        \cache[7][2][TAG][6] ), .ZN(n744) );
  NAND4_X1 U951 ( .A1(n747), .A2(n746), .A3(n745), .A4(n744), .ZN(n749) );
  AOI22_X1 U952 ( .A1(pc_fetch[9]), .A2(n751), .B1(n749), .B2(n750), .ZN(n748)
         );
  OAI221_X1 U953 ( .B1(pc_fetch[9]), .B2(n751), .C1(n750), .C2(n749), .A(n748), 
        .ZN(n806) );
  AOI22_X1 U954 ( .A1(n234), .A2(\cache[0][2][TAG][7] ), .B1(n36), .B2(
        \cache[1][2][TAG][7] ), .ZN(n755) );
  AOI22_X1 U955 ( .A1(n55), .A2(\cache[2][2][TAG][7] ), .B1(n37), .B2(
        \cache[3][2][TAG][7] ), .ZN(n754) );
  AOI22_X1 U956 ( .A1(n56), .A2(\cache[4][2][TAG][7] ), .B1(n38), .B2(
        \cache[5][2][TAG][7] ), .ZN(n753) );
  AOI22_X1 U957 ( .A1(n40), .A2(\cache[6][2][TAG][7] ), .B1(n39), .B2(
        \cache[7][2][TAG][7] ), .ZN(n752) );
  AND4_X1 U958 ( .A1(n755), .A2(n754), .A3(n753), .A4(n752), .ZN(n762) );
  AOI22_X1 U959 ( .A1(n234), .A2(\cache[0][2][TAG][5] ), .B1(n36), .B2(
        \cache[1][2][TAG][5] ), .ZN(n759) );
  AOI22_X1 U960 ( .A1(n239), .A2(\cache[2][2][TAG][5] ), .B1(n37), .B2(
        \cache[3][2][TAG][5] ), .ZN(n758) );
  AOI22_X1 U961 ( .A1(n243), .A2(\cache[4][2][TAG][5] ), .B1(n38), .B2(
        \cache[5][2][TAG][5] ), .ZN(n757) );
  AOI22_X1 U962 ( .A1(n40), .A2(\cache[6][2][TAG][5] ), .B1(n39), .B2(
        \cache[7][2][TAG][5] ), .ZN(n756) );
  NAND4_X1 U963 ( .A1(n759), .A2(n758), .A3(n757), .A4(n756), .ZN(n761) );
  AOI22_X1 U964 ( .A1(pc_fetch[12]), .A2(n762), .B1(n761), .B2(n65), .ZN(n760)
         );
  OAI221_X1 U965 ( .B1(pc_fetch[12]), .B2(n762), .C1(n65), .C2(n761), .A(n760), 
        .ZN(n805) );
  AOI22_X1 U966 ( .A1(n234), .A2(\cache[0][2][TAG][1] ), .B1(n36), .B2(
        \cache[1][2][TAG][1] ), .ZN(n766) );
  AOI22_X1 U967 ( .A1(n1571), .A2(\cache[2][2][TAG][1] ), .B1(n37), .B2(
        \cache[3][2][TAG][1] ), .ZN(n765) );
  AOI22_X1 U968 ( .A1(n1573), .A2(\cache[4][2][TAG][1] ), .B1(n38), .B2(
        \cache[5][2][TAG][1] ), .ZN(n764) );
  AOI22_X1 U969 ( .A1(n40), .A2(\cache[6][2][TAG][1] ), .B1(n39), .B2(
        \cache[7][2][TAG][1] ), .ZN(n763) );
  AND4_X1 U970 ( .A1(n766), .A2(n765), .A3(n764), .A4(n763), .ZN(n773) );
  AOI22_X1 U971 ( .A1(n234), .A2(\cache[0][2][TAG][3] ), .B1(n36), .B2(
        \cache[1][2][TAG][3] ), .ZN(n770) );
  AOI22_X1 U972 ( .A1(n239), .A2(\cache[2][2][TAG][3] ), .B1(n37), .B2(
        \cache[3][2][TAG][3] ), .ZN(n769) );
  AOI22_X1 U973 ( .A1(n243), .A2(\cache[4][2][TAG][3] ), .B1(n38), .B2(
        \cache[5][2][TAG][3] ), .ZN(n768) );
  AOI22_X1 U974 ( .A1(n40), .A2(\cache[6][2][TAG][3] ), .B1(n39), .B2(
        \cache[7][2][TAG][3] ), .ZN(n767) );
  NAND4_X1 U975 ( .A1(n770), .A2(n769), .A3(n768), .A4(n767), .ZN(n772) );
  AOI22_X1 U976 ( .A1(pc_fetch[6]), .A2(n773), .B1(n772), .B2(n66), .ZN(n771)
         );
  OAI221_X1 U977 ( .B1(pc_fetch[6]), .B2(n773), .C1(n66), .C2(n772), .A(n771), 
        .ZN(n804) );
  AOI22_X1 U978 ( .A1(\cache[0][2][YOUTH][2] ), .A2(n57), .B1(
        \cache[1][2][YOUTH][2] ), .B2(n36), .ZN(n777) );
  AOI22_X1 U979 ( .A1(\cache[3][2][YOUTH][2] ), .A2(n37), .B1(
        \cache[2][2][YOUTH][2] ), .B2(n1571), .ZN(n776) );
  AOI22_X1 U980 ( .A1(\cache[5][2][YOUTH][2] ), .A2(n38), .B1(
        \cache[4][2][YOUTH][2] ), .B2(n1573), .ZN(n775) );
  AOI22_X1 U981 ( .A1(\cache[7][2][YOUTH][2] ), .A2(n39), .B1(
        \cache[6][2][YOUTH][2] ), .B2(n40), .ZN(n774) );
  NAND4_X1 U982 ( .A1(n777), .A2(n776), .A3(n775), .A4(n774), .ZN(n788) );
  AOI22_X1 U983 ( .A1(\cache[0][2][YOUTH][0] ), .A2(n57), .B1(
        \cache[1][2][YOUTH][0] ), .B2(n36), .ZN(n781) );
  AOI22_X1 U984 ( .A1(\cache[3][2][YOUTH][0] ), .A2(n37), .B1(
        \cache[2][2][YOUTH][0] ), .B2(n1571), .ZN(n780) );
  AOI22_X1 U985 ( .A1(\cache[5][2][YOUTH][0] ), .A2(n38), .B1(
        \cache[4][2][YOUTH][0] ), .B2(n1573), .ZN(n779) );
  AOI22_X1 U986 ( .A1(\cache[7][2][YOUTH][0] ), .A2(n39), .B1(
        \cache[6][2][YOUTH][0] ), .B2(n40), .ZN(n778) );
  NAND4_X1 U987 ( .A1(n781), .A2(n780), .A3(n779), .A4(n778), .ZN(n787) );
  AOI22_X1 U988 ( .A1(\cache[0][2][YOUTH][1] ), .A2(n57), .B1(
        \cache[1][2][YOUTH][1] ), .B2(n36), .ZN(n785) );
  AOI22_X1 U989 ( .A1(\cache[3][2][YOUTH][1] ), .A2(n37), .B1(
        \cache[2][2][YOUTH][1] ), .B2(n1571), .ZN(n784) );
  AOI22_X1 U990 ( .A1(\cache[5][2][YOUTH][1] ), .A2(n38), .B1(
        \cache[4][2][YOUTH][1] ), .B2(n1573), .ZN(n783) );
  AOI22_X1 U991 ( .A1(\cache[7][2][YOUTH][1] ), .A2(n39), .B1(
        \cache[6][2][YOUTH][1] ), .B2(n40), .ZN(n782) );
  NAND4_X1 U992 ( .A1(n785), .A2(n784), .A3(n783), .A4(n782), .ZN(n786) );
  NAND3_X1 U993 ( .A1(n788), .A2(n787), .A3(n786), .ZN(n802) );
  AOI22_X1 U994 ( .A1(n57), .A2(\cache[0][2][TAG][0] ), .B1(n36), .B2(
        \cache[1][2][TAG][0] ), .ZN(n792) );
  AOI22_X1 U995 ( .A1(n55), .A2(\cache[2][2][TAG][0] ), .B1(n37), .B2(
        \cache[3][2][TAG][0] ), .ZN(n791) );
  AOI22_X1 U996 ( .A1(n56), .A2(\cache[4][2][TAG][0] ), .B1(n38), .B2(
        \cache[5][2][TAG][0] ), .ZN(n790) );
  AOI22_X1 U997 ( .A1(n40), .A2(\cache[6][2][TAG][0] ), .B1(n39), .B2(
        \cache[7][2][TAG][0] ), .ZN(n789) );
  NAND4_X1 U998 ( .A1(n792), .A2(n791), .A3(n790), .A4(n789), .ZN(n800) );
  AOI22_X1 U999 ( .A1(n57), .A2(\cache[0][2][TAG][2] ), .B1(n36), .B2(
        \cache[1][2][TAG][2] ), .ZN(n796) );
  AOI22_X1 U1000 ( .A1(n55), .A2(\cache[2][2][TAG][2] ), .B1(n37), .B2(
        \cache[3][2][TAG][2] ), .ZN(n795) );
  AOI22_X1 U1001 ( .A1(n56), .A2(\cache[4][2][TAG][2] ), .B1(n38), .B2(
        \cache[5][2][TAG][2] ), .ZN(n794) );
  AOI22_X1 U1002 ( .A1(n40), .A2(\cache[6][2][TAG][2] ), .B1(n39), .B2(
        \cache[7][2][TAG][2] ), .ZN(n793) );
  AND4_X1 U1003 ( .A1(n796), .A2(n795), .A3(n794), .A4(n793), .ZN(n798) );
  OAI22_X1 U1004 ( .A1(n799), .A2(n800), .B1(pc_fetch[7]), .B2(n798), .ZN(n797) );
  AOI221_X1 U1005 ( .B1(n800), .B2(n799), .C1(pc_fetch[7]), .C2(n798), .A(n797), .ZN(n801) );
  NAND2_X1 U1006 ( .A1(n802), .A2(n801), .ZN(n803) );
  NOR4_X1 U1007 ( .A1(n806), .A2(n805), .A3(n804), .A4(n803), .ZN(n809) );
  AND2_X1 U1008 ( .A1(n884), .A2(n809), .ZN(n895) );
  OAI21_X1 U1009 ( .B1(n807), .B2(n895), .A(n882), .ZN(\hit_index[0] ) );
  INV_X1 U1010 ( .A(n807), .ZN(n886) );
  NAND2_X1 U1011 ( .A1(n884), .A2(n886), .ZN(n808) );
  NAND2_X1 U1012 ( .A1(n882), .A2(n808), .ZN(\hit_index[1] ) );
  NOR2_X1 U1013 ( .A1(n809), .A2(n808), .ZN(n900) );
  AOI22_X1 U1014 ( .A1(n57), .A2(\cache[0][3][TAG][3] ), .B1(n36), .B2(
        \cache[1][3][TAG][3] ), .ZN(n813) );
  AOI22_X1 U1015 ( .A1(n55), .A2(\cache[2][3][TAG][3] ), .B1(n37), .B2(
        \cache[3][3][TAG][3] ), .ZN(n812) );
  AOI22_X1 U1016 ( .A1(n56), .A2(\cache[4][3][TAG][3] ), .B1(n38), .B2(
        \cache[5][3][TAG][3] ), .ZN(n811) );
  AOI22_X1 U1017 ( .A1(n40), .A2(\cache[6][3][TAG][3] ), .B1(n39), .B2(
        \cache[7][3][TAG][3] ), .ZN(n810) );
  NAND4_X1 U1018 ( .A1(n813), .A2(n812), .A3(n811), .A4(n810), .ZN(n820) );
  AOI22_X1 U1019 ( .A1(n236), .A2(\cache[0][3][TAG][2] ), .B1(n36), .B2(
        \cache[1][3][TAG][2] ), .ZN(n817) );
  AOI22_X1 U1020 ( .A1(n55), .A2(\cache[2][3][TAG][2] ), .B1(n37), .B2(
        \cache[3][3][TAG][2] ), .ZN(n816) );
  AOI22_X1 U1021 ( .A1(n56), .A2(\cache[4][3][TAG][2] ), .B1(n38), .B2(
        \cache[5][3][TAG][2] ), .ZN(n815) );
  AOI22_X1 U1022 ( .A1(n40), .A2(\cache[6][3][TAG][2] ), .B1(n39), .B2(
        \cache[7][3][TAG][2] ), .ZN(n814) );
  AND4_X1 U1023 ( .A1(n817), .A2(n816), .A3(n815), .A4(n814), .ZN(n819) );
  OAI22_X1 U1024 ( .A1(n66), .A2(n820), .B1(n819), .B2(pc_fetch[7]), .ZN(n818)
         );
  AOI221_X1 U1025 ( .B1(n820), .B2(n66), .C1(n819), .C2(pc_fetch[7]), .A(n818), 
        .ZN(n875) );
  AOI22_X1 U1026 ( .A1(n236), .A2(\cache[0][3][TAG][1] ), .B1(n36), .B2(
        \cache[1][3][TAG][1] ), .ZN(n824) );
  AOI22_X1 U1027 ( .A1(n55), .A2(\cache[2][3][TAG][1] ), .B1(n37), .B2(
        \cache[3][3][TAG][1] ), .ZN(n823) );
  AOI22_X1 U1028 ( .A1(n56), .A2(\cache[4][3][TAG][1] ), .B1(n38), .B2(
        \cache[5][3][TAG][1] ), .ZN(n822) );
  AOI22_X1 U1029 ( .A1(n40), .A2(\cache[6][3][TAG][1] ), .B1(n39), .B2(
        \cache[7][3][TAG][1] ), .ZN(n821) );
  NAND4_X1 U1030 ( .A1(n824), .A2(n823), .A3(n822), .A4(n821), .ZN(n831) );
  AOI22_X1 U1031 ( .A1(n236), .A2(\cache[0][3][TAG][0] ), .B1(n36), .B2(
        \cache[1][3][TAG][0] ), .ZN(n828) );
  AOI22_X1 U1032 ( .A1(n55), .A2(\cache[2][3][TAG][0] ), .B1(n37), .B2(
        \cache[3][3][TAG][0] ), .ZN(n827) );
  AOI22_X1 U1033 ( .A1(n56), .A2(\cache[4][3][TAG][0] ), .B1(n38), .B2(
        \cache[5][3][TAG][0] ), .ZN(n826) );
  AOI22_X1 U1034 ( .A1(n40), .A2(\cache[6][3][TAG][0] ), .B1(n39), .B2(
        \cache[7][3][TAG][0] ), .ZN(n825) );
  AND4_X1 U1035 ( .A1(n828), .A2(n827), .A3(n826), .A4(n825), .ZN(n830) );
  OAI22_X1 U1036 ( .A1(n67), .A2(n831), .B1(pc_fetch[5]), .B2(n830), .ZN(n829)
         );
  AOI221_X1 U1037 ( .B1(n831), .B2(n67), .C1(pc_fetch[5]), .C2(n830), .A(n829), 
        .ZN(n874) );
  AOI22_X1 U1038 ( .A1(n234), .A2(\cache[0][3][TAG][4] ), .B1(n36), .B2(
        \cache[1][3][TAG][4] ), .ZN(n835) );
  AOI22_X1 U1039 ( .A1(n55), .A2(\cache[2][3][TAG][4] ), .B1(n37), .B2(
        \cache[3][3][TAG][4] ), .ZN(n834) );
  AOI22_X1 U1040 ( .A1(n56), .A2(\cache[4][3][TAG][4] ), .B1(n38), .B2(
        \cache[5][3][TAG][4] ), .ZN(n833) );
  AOI22_X1 U1041 ( .A1(n40), .A2(\cache[6][3][TAG][4] ), .B1(n39), .B2(
        \cache[7][3][TAG][4] ), .ZN(n832) );
  AND4_X1 U1042 ( .A1(n835), .A2(n834), .A3(n833), .A4(n832), .ZN(n842) );
  AOI22_X1 U1043 ( .A1(n57), .A2(\cache[0][3][TAG][5] ), .B1(n36), .B2(
        \cache[1][3][TAG][5] ), .ZN(n839) );
  AOI22_X1 U1044 ( .A1(n55), .A2(\cache[2][3][TAG][5] ), .B1(n37), .B2(
        \cache[3][3][TAG][5] ), .ZN(n838) );
  AOI22_X1 U1045 ( .A1(n56), .A2(\cache[4][3][TAG][5] ), .B1(n38), .B2(
        \cache[5][3][TAG][5] ), .ZN(n837) );
  AOI22_X1 U1046 ( .A1(n40), .A2(\cache[6][3][TAG][5] ), .B1(n39), .B2(
        \cache[7][3][TAG][5] ), .ZN(n836) );
  NAND4_X1 U1047 ( .A1(n839), .A2(n838), .A3(n837), .A4(n836), .ZN(n841) );
  AOI22_X1 U1048 ( .A1(pc_fetch[9]), .A2(n842), .B1(n841), .B2(n65), .ZN(n840)
         );
  OAI221_X1 U1049 ( .B1(pc_fetch[9]), .B2(n842), .C1(n65), .C2(n841), .A(n840), 
        .ZN(n856) );
  AOI22_X1 U1050 ( .A1(n234), .A2(\cache[0][3][TAG][6] ), .B1(n36), .B2(
        \cache[1][3][TAG][6] ), .ZN(n846) );
  AOI22_X1 U1051 ( .A1(n55), .A2(\cache[2][3][TAG][6] ), .B1(n37), .B2(
        \cache[3][3][TAG][6] ), .ZN(n845) );
  AOI22_X1 U1052 ( .A1(n56), .A2(\cache[4][3][TAG][6] ), .B1(n38), .B2(
        \cache[5][3][TAG][6] ), .ZN(n844) );
  AOI22_X1 U1053 ( .A1(n40), .A2(\cache[6][3][TAG][6] ), .B1(n39), .B2(
        \cache[7][3][TAG][6] ), .ZN(n843) );
  AND4_X1 U1054 ( .A1(n846), .A2(n845), .A3(n844), .A4(n843), .ZN(n854) );
  AOI22_X1 U1055 ( .A1(n234), .A2(\cache[0][3][TAG][7] ), .B1(n36), .B2(
        \cache[1][3][TAG][7] ), .ZN(n851) );
  AOI22_X1 U1056 ( .A1(n55), .A2(\cache[2][3][TAG][7] ), .B1(n37), .B2(
        \cache[3][3][TAG][7] ), .ZN(n850) );
  AOI22_X1 U1057 ( .A1(n56), .A2(\cache[4][3][TAG][7] ), .B1(n38), .B2(
        \cache[5][3][TAG][7] ), .ZN(n848) );
  AOI22_X1 U1058 ( .A1(n40), .A2(\cache[6][3][TAG][7] ), .B1(n39), .B2(
        \cache[7][3][TAG][7] ), .ZN(n847) );
  NAND4_X1 U1059 ( .A1(n851), .A2(n850), .A3(n848), .A4(n847), .ZN(n853) );
  AOI22_X1 U1060 ( .A1(pc_fetch[11]), .A2(n854), .B1(n853), .B2(n64), .ZN(n852) );
  OAI221_X1 U1061 ( .B1(pc_fetch[11]), .B2(n854), .C1(n64), .C2(n853), .A(n852), .ZN(n855) );
  NOR2_X1 U1062 ( .A1(n856), .A2(n855), .ZN(n873) );
  AOI22_X1 U1063 ( .A1(\cache[0][3][YOUTH][2] ), .A2(n57), .B1(
        \cache[1][3][YOUTH][2] ), .B2(n36), .ZN(n860) );
  AOI22_X1 U1064 ( .A1(\cache[3][3][YOUTH][2] ), .A2(n37), .B1(
        \cache[2][3][YOUTH][2] ), .B2(n239), .ZN(n859) );
  AOI22_X1 U1065 ( .A1(\cache[5][3][YOUTH][2] ), .A2(n38), .B1(
        \cache[4][3][YOUTH][2] ), .B2(n243), .ZN(n858) );
  AOI22_X1 U1066 ( .A1(\cache[7][3][YOUTH][2] ), .A2(n39), .B1(
        \cache[6][3][YOUTH][2] ), .B2(n40), .ZN(n857) );
  NAND4_X1 U1067 ( .A1(n860), .A2(n859), .A3(n858), .A4(n857), .ZN(n871) );
  AOI22_X1 U1068 ( .A1(\cache[0][3][YOUTH][0] ), .A2(n57), .B1(
        \cache[1][3][YOUTH][0] ), .B2(n36), .ZN(n864) );
  AOI22_X1 U1069 ( .A1(\cache[3][3][YOUTH][0] ), .A2(n37), .B1(
        \cache[2][3][YOUTH][0] ), .B2(n239), .ZN(n863) );
  AOI22_X1 U1070 ( .A1(\cache[5][3][YOUTH][0] ), .A2(n38), .B1(
        \cache[4][3][YOUTH][0] ), .B2(n243), .ZN(n862) );
  AOI22_X1 U1071 ( .A1(\cache[7][3][YOUTH][0] ), .A2(n39), .B1(
        \cache[6][3][YOUTH][0] ), .B2(n40), .ZN(n861) );
  NAND4_X1 U1072 ( .A1(n864), .A2(n863), .A3(n862), .A4(n861), .ZN(n870) );
  AOI22_X1 U1073 ( .A1(\cache[0][3][YOUTH][1] ), .A2(n236), .B1(
        \cache[1][3][YOUTH][1] ), .B2(n36), .ZN(n868) );
  AOI22_X1 U1074 ( .A1(\cache[3][3][YOUTH][1] ), .A2(n37), .B1(
        \cache[2][3][YOUTH][1] ), .B2(n240), .ZN(n867) );
  AOI22_X1 U1075 ( .A1(\cache[5][3][YOUTH][1] ), .A2(n38), .B1(
        \cache[4][3][YOUTH][1] ), .B2(n244), .ZN(n866) );
  AOI22_X1 U1076 ( .A1(\cache[7][3][YOUTH][1] ), .A2(n39), .B1(
        \cache[6][3][YOUTH][1] ), .B2(n40), .ZN(n865) );
  NAND4_X1 U1077 ( .A1(n868), .A2(n867), .A3(n866), .A4(n865), .ZN(n869) );
  NAND3_X1 U1078 ( .A1(n871), .A2(n870), .A3(n869), .ZN(n872) );
  NAND4_X1 U1079 ( .A1(n875), .A2(n874), .A3(n873), .A4(n872), .ZN(n901) );
  NAND2_X1 U1080 ( .A1(n900), .A2(n901), .ZN(n883) );
  NAND2_X1 U1081 ( .A1(n882), .A2(n883), .ZN(\hit_index[2] ) );
  AOI21_X1 U1082 ( .B1(n906), .B2(n883), .A(n201), .ZN(n1118) );
  NAND2_X1 U1083 ( .A1(n1118), .A2(pc_in[0]), .ZN(n876) );
  OAI21_X1 U1084 ( .B1(n877), .B2(n88), .A(n876), .ZN(pc_out[0]) );
  INV_X1 U1085 ( .A(pc_out[0]), .ZN(n849) );
  AOI22_X1 U1086 ( .A1(n57), .A2(\cache[0][1][DATA][8] ), .B1(n36), .B2(
        \cache[1][1][DATA][8] ), .ZN(n881) );
  AOI22_X1 U1087 ( .A1(n240), .A2(\cache[2][1][DATA][8] ), .B1(n37), .B2(
        \cache[3][1][DATA][8] ), .ZN(n880) );
  AOI22_X1 U1088 ( .A1(n244), .A2(\cache[4][1][DATA][8] ), .B1(n38), .B2(
        \cache[5][1][DATA][8] ), .ZN(n879) );
  AOI22_X1 U1089 ( .A1(n40), .A2(\cache[6][1][DATA][8] ), .B1(n39), .B2(
        \cache[7][1][DATA][8] ), .ZN(n878) );
  AND4_X1 U1090 ( .A1(n881), .A2(n880), .A3(n879), .A4(n878), .ZN(n910) );
  AOI22_X1 U1091 ( .A1(n57), .A2(\cache[0][0][DATA][8] ), .B1(n36), .B2(
        \cache[1][0][DATA][8] ), .ZN(n890) );
  AOI22_X1 U1092 ( .A1(n240), .A2(\cache[2][0][DATA][8] ), .B1(n37), .B2(
        \cache[3][0][DATA][8] ), .ZN(n889) );
  AOI22_X1 U1093 ( .A1(n244), .A2(\cache[4][0][DATA][8] ), .B1(n38), .B2(
        \cache[5][0][DATA][8] ), .ZN(n888) );
  AOI22_X1 U1094 ( .A1(n40), .A2(\cache[6][0][DATA][8] ), .B1(n39), .B2(
        \cache[7][0][DATA][8] ), .ZN(n887) );
  NAND4_X1 U1095 ( .A1(n890), .A2(n889), .A3(n888), .A4(n887), .ZN(n899) );
  AOI22_X1 U1096 ( .A1(n1569), .A2(\cache[0][2][DATA][8] ), .B1(n36), .B2(
        \cache[1][2][DATA][8] ), .ZN(n894) );
  AOI22_X1 U1097 ( .A1(n240), .A2(\cache[2][2][DATA][8] ), .B1(n37), .B2(
        \cache[3][2][DATA][8] ), .ZN(n893) );
  AOI22_X1 U1098 ( .A1(n244), .A2(\cache[4][2][DATA][8] ), .B1(n38), .B2(
        \cache[5][2][DATA][8] ), .ZN(n892) );
  AOI22_X1 U1099 ( .A1(n40), .A2(\cache[6][2][DATA][8] ), .B1(n39), .B2(
        \cache[7][2][DATA][8] ), .ZN(n891) );
  AND4_X1 U1100 ( .A1(n894), .A2(n893), .A3(n892), .A4(n891), .ZN(n897) );
  NAND2_X1 U1101 ( .A1(n896), .A2(n895), .ZN(n1563) );
  OAI22_X1 U1102 ( .A1(n897), .A2(n227), .B1(n271), .B2(n87), .ZN(n898) );
  AOI21_X1 U1103 ( .B1(n229), .B2(n899), .A(n898), .ZN(n909) );
  AOI22_X1 U1104 ( .A1(n57), .A2(\cache[0][3][DATA][8] ), .B1(n36), .B2(
        \cache[1][3][DATA][8] ), .ZN(n905) );
  AOI22_X1 U1105 ( .A1(n240), .A2(\cache[2][3][DATA][8] ), .B1(n37), .B2(
        \cache[3][3][DATA][8] ), .ZN(n904) );
  AOI22_X1 U1106 ( .A1(n244), .A2(\cache[4][3][DATA][8] ), .B1(n38), .B2(
        \cache[5][3][DATA][8] ), .ZN(n903) );
  AOI22_X1 U1107 ( .A1(n40), .A2(\cache[6][3][DATA][8] ), .B1(n39), .B2(
        \cache[7][3][DATA][8] ), .ZN(n902) );
  NAND4_X1 U1108 ( .A1(n905), .A2(n904), .A3(n903), .A4(n902), .ZN(n907) );
  AOI22_X1 U1109 ( .A1(n249), .A2(n907), .B1(pc_in[10]), .B2(n93), .ZN(n908)
         );
  OAI211_X1 U1110 ( .C1(n910), .C2(n1584), .A(n909), .B(n908), .ZN(pc_out[10])
         );
  AOI22_X1 U1111 ( .A1(n57), .A2(\cache[0][1][DATA][9] ), .B1(n36), .B2(
        \cache[1][1][DATA][9] ), .ZN(n914) );
  AOI22_X1 U1112 ( .A1(n240), .A2(\cache[2][1][DATA][9] ), .B1(n37), .B2(
        \cache[3][1][DATA][9] ), .ZN(n913) );
  AOI22_X1 U1113 ( .A1(n244), .A2(\cache[4][1][DATA][9] ), .B1(n38), .B2(
        \cache[5][1][DATA][9] ), .ZN(n912) );
  AOI22_X1 U1114 ( .A1(n40), .A2(\cache[6][1][DATA][9] ), .B1(n39), .B2(
        \cache[7][1][DATA][9] ), .ZN(n911) );
  AND4_X1 U1115 ( .A1(n914), .A2(n913), .A3(n912), .A4(n911), .ZN(n933) );
  AOI22_X1 U1116 ( .A1(n235), .A2(\cache[0][0][DATA][9] ), .B1(n36), .B2(
        \cache[1][0][DATA][9] ), .ZN(n918) );
  AOI22_X1 U1117 ( .A1(n240), .A2(\cache[2][0][DATA][9] ), .B1(n37), .B2(
        \cache[3][0][DATA][9] ), .ZN(n917) );
  AOI22_X1 U1118 ( .A1(n244), .A2(\cache[4][0][DATA][9] ), .B1(n38), .B2(
        \cache[5][0][DATA][9] ), .ZN(n916) );
  AOI22_X1 U1119 ( .A1(n40), .A2(\cache[6][0][DATA][9] ), .B1(n39), .B2(
        \cache[7][0][DATA][9] ), .ZN(n915) );
  NAND4_X1 U1120 ( .A1(n918), .A2(n917), .A3(n916), .A4(n915), .ZN(n925) );
  AOI22_X1 U1121 ( .A1(n1569), .A2(\cache[0][2][DATA][9] ), .B1(n36), .B2(
        \cache[1][2][DATA][9] ), .ZN(n922) );
  AOI22_X1 U1122 ( .A1(n240), .A2(\cache[2][2][DATA][9] ), .B1(n37), .B2(
        \cache[3][2][DATA][9] ), .ZN(n921) );
  AOI22_X1 U1123 ( .A1(n244), .A2(\cache[4][2][DATA][9] ), .B1(n38), .B2(
        \cache[5][2][DATA][9] ), .ZN(n920) );
  AOI22_X1 U1124 ( .A1(n40), .A2(\cache[6][2][DATA][9] ), .B1(n39), .B2(
        \cache[7][2][DATA][9] ), .ZN(n919) );
  AND4_X1 U1125 ( .A1(n922), .A2(n921), .A3(n920), .A4(n919), .ZN(n923) );
  OAI22_X1 U1126 ( .A1(n923), .A2(n228), .B1(n272), .B2(n87), .ZN(n924) );
  AOI21_X1 U1127 ( .B1(n25), .B2(n925), .A(n924), .ZN(n932) );
  AOI22_X1 U1128 ( .A1(n235), .A2(\cache[0][3][DATA][9] ), .B1(n36), .B2(
        \cache[1][3][DATA][9] ), .ZN(n929) );
  AOI22_X1 U1129 ( .A1(n240), .A2(\cache[2][3][DATA][9] ), .B1(n37), .B2(
        \cache[3][3][DATA][9] ), .ZN(n928) );
  AOI22_X1 U1130 ( .A1(n244), .A2(\cache[4][3][DATA][9] ), .B1(n38), .B2(
        \cache[5][3][DATA][9] ), .ZN(n927) );
  AOI22_X1 U1131 ( .A1(n40), .A2(\cache[6][3][DATA][9] ), .B1(n39), .B2(
        \cache[7][3][DATA][9] ), .ZN(n926) );
  NAND4_X1 U1132 ( .A1(n929), .A2(n928), .A3(n927), .A4(n926), .ZN(n930) );
  AOI22_X1 U1133 ( .A1(n248), .A2(n930), .B1(pc_in[11]), .B2(n93), .ZN(n931)
         );
  OAI211_X1 U1134 ( .C1(n933), .C2(n1584), .A(n932), .B(n931), .ZN(pc_out[11])
         );
  AOI22_X1 U1135 ( .A1(n57), .A2(\cache[0][1][DATA][10] ), .B1(n36), .B2(
        \cache[1][1][DATA][10] ), .ZN(n937) );
  AOI22_X1 U1136 ( .A1(n240), .A2(\cache[2][1][DATA][10] ), .B1(n37), .B2(
        \cache[3][1][DATA][10] ), .ZN(n936) );
  AOI22_X1 U1137 ( .A1(n244), .A2(\cache[4][1][DATA][10] ), .B1(n38), .B2(
        \cache[5][1][DATA][10] ), .ZN(n935) );
  AOI22_X1 U1138 ( .A1(n40), .A2(\cache[6][1][DATA][10] ), .B1(n39), .B2(
        \cache[7][1][DATA][10] ), .ZN(n934) );
  AND4_X1 U1139 ( .A1(n937), .A2(n936), .A3(n935), .A4(n934), .ZN(n956) );
  AOI22_X1 U1140 ( .A1(n57), .A2(\cache[0][0][DATA][10] ), .B1(n36), .B2(
        \cache[1][0][DATA][10] ), .ZN(n941) );
  AOI22_X1 U1141 ( .A1(n240), .A2(\cache[2][0][DATA][10] ), .B1(n37), .B2(
        \cache[3][0][DATA][10] ), .ZN(n940) );
  AOI22_X1 U1142 ( .A1(n244), .A2(\cache[4][0][DATA][10] ), .B1(n38), .B2(
        \cache[5][0][DATA][10] ), .ZN(n939) );
  AOI22_X1 U1143 ( .A1(n40), .A2(\cache[6][0][DATA][10] ), .B1(n39), .B2(
        \cache[7][0][DATA][10] ), .ZN(n938) );
  NAND4_X1 U1144 ( .A1(n941), .A2(n940), .A3(n939), .A4(n938), .ZN(n948) );
  AOI22_X1 U1145 ( .A1(n1569), .A2(\cache[0][2][DATA][10] ), .B1(n36), .B2(
        \cache[1][2][DATA][10] ), .ZN(n945) );
  AOI22_X1 U1146 ( .A1(n240), .A2(\cache[2][2][DATA][10] ), .B1(n37), .B2(
        \cache[3][2][DATA][10] ), .ZN(n944) );
  AOI22_X1 U1147 ( .A1(n244), .A2(\cache[4][2][DATA][10] ), .B1(n38), .B2(
        \cache[5][2][DATA][10] ), .ZN(n943) );
  AOI22_X1 U1148 ( .A1(n40), .A2(\cache[6][2][DATA][10] ), .B1(n39), .B2(
        \cache[7][2][DATA][10] ), .ZN(n942) );
  AND4_X1 U1149 ( .A1(n945), .A2(n944), .A3(n943), .A4(n942), .ZN(n946) );
  OAI22_X1 U1150 ( .A1(n946), .A2(n227), .B1(n273), .B2(n87), .ZN(n947) );
  AOI21_X1 U1151 ( .B1(n230), .B2(n948), .A(n947), .ZN(n955) );
  AOI22_X1 U1152 ( .A1(n57), .A2(\cache[0][3][DATA][10] ), .B1(n36), .B2(
        \cache[1][3][DATA][10] ), .ZN(n952) );
  AOI22_X1 U1153 ( .A1(n240), .A2(\cache[2][3][DATA][10] ), .B1(n37), .B2(
        \cache[3][3][DATA][10] ), .ZN(n951) );
  AOI22_X1 U1154 ( .A1(n244), .A2(\cache[4][3][DATA][10] ), .B1(n38), .B2(
        \cache[5][3][DATA][10] ), .ZN(n950) );
  AOI22_X1 U1155 ( .A1(n40), .A2(\cache[6][3][DATA][10] ), .B1(n39), .B2(
        \cache[7][3][DATA][10] ), .ZN(n949) );
  NAND4_X1 U1156 ( .A1(n952), .A2(n951), .A3(n950), .A4(n949), .ZN(n953) );
  AOI22_X1 U1157 ( .A1(n248), .A2(n953), .B1(pc_in[12]), .B2(n93), .ZN(n954)
         );
  OAI211_X1 U1158 ( .C1(n956), .C2(n1584), .A(n955), .B(n954), .ZN(pc_out[12])
         );
  AOI22_X1 U1159 ( .A1(n235), .A2(\cache[0][1][DATA][11] ), .B1(n232), .B2(
        \cache[1][1][DATA][11] ), .ZN(n960) );
  AOI22_X1 U1160 ( .A1(n55), .A2(\cache[2][1][DATA][11] ), .B1(n37), .B2(
        \cache[3][1][DATA][11] ), .ZN(n959) );
  AOI22_X1 U1161 ( .A1(n56), .A2(\cache[4][1][DATA][11] ), .B1(n38), .B2(
        \cache[5][1][DATA][11] ), .ZN(n958) );
  AOI22_X1 U1162 ( .A1(n40), .A2(\cache[6][1][DATA][11] ), .B1(n246), .B2(
        \cache[7][1][DATA][11] ), .ZN(n957) );
  AND4_X1 U1163 ( .A1(n960), .A2(n959), .A3(n958), .A4(n957), .ZN(n979) );
  AOI22_X1 U1164 ( .A1(n236), .A2(\cache[0][0][DATA][11] ), .B1(n36), .B2(
        \cache[1][0][DATA][11] ), .ZN(n964) );
  AOI22_X1 U1165 ( .A1(n240), .A2(\cache[2][0][DATA][11] ), .B1(n37), .B2(
        \cache[3][0][DATA][11] ), .ZN(n963) );
  AOI22_X1 U1166 ( .A1(n56), .A2(\cache[4][0][DATA][11] ), .B1(n38), .B2(
        \cache[5][0][DATA][11] ), .ZN(n962) );
  AOI22_X1 U1167 ( .A1(n40), .A2(\cache[6][0][DATA][11] ), .B1(n246), .B2(
        \cache[7][0][DATA][11] ), .ZN(n961) );
  NAND4_X1 U1168 ( .A1(n964), .A2(n963), .A3(n962), .A4(n961), .ZN(n971) );
  AOI22_X1 U1169 ( .A1(n235), .A2(\cache[0][2][DATA][11] ), .B1(n36), .B2(
        \cache[1][2][DATA][11] ), .ZN(n968) );
  AOI22_X1 U1170 ( .A1(n240), .A2(\cache[2][2][DATA][11] ), .B1(n37), .B2(
        \cache[3][2][DATA][11] ), .ZN(n967) );
  AOI22_X1 U1171 ( .A1(n244), .A2(\cache[4][2][DATA][11] ), .B1(n38), .B2(
        \cache[5][2][DATA][11] ), .ZN(n966) );
  AOI22_X1 U1172 ( .A1(n40), .A2(\cache[6][2][DATA][11] ), .B1(n39), .B2(
        \cache[7][2][DATA][11] ), .ZN(n965) );
  AND4_X1 U1173 ( .A1(n968), .A2(n967), .A3(n966), .A4(n965), .ZN(n969) );
  OAI22_X1 U1174 ( .A1(n969), .A2(n228), .B1(n274), .B2(n87), .ZN(n970) );
  AOI21_X1 U1175 ( .B1(n230), .B2(n971), .A(n970), .ZN(n978) );
  AOI22_X1 U1176 ( .A1(n233), .A2(\cache[0][3][DATA][11] ), .B1(n232), .B2(
        \cache[1][3][DATA][11] ), .ZN(n975) );
  AOI22_X1 U1177 ( .A1(n240), .A2(\cache[2][3][DATA][11] ), .B1(n237), .B2(
        \cache[3][3][DATA][11] ), .ZN(n974) );
  AOI22_X1 U1178 ( .A1(n244), .A2(\cache[4][3][DATA][11] ), .B1(n241), .B2(
        \cache[5][3][DATA][11] ), .ZN(n973) );
  AOI22_X1 U1179 ( .A1(n40), .A2(\cache[6][3][DATA][11] ), .B1(n39), .B2(
        \cache[7][3][DATA][11] ), .ZN(n972) );
  NAND4_X1 U1180 ( .A1(n975), .A2(n974), .A3(n973), .A4(n972), .ZN(n976) );
  AOI22_X1 U1181 ( .A1(n249), .A2(n976), .B1(pc_in[13]), .B2(n93), .ZN(n977)
         );
  OAI211_X1 U1182 ( .C1(n979), .C2(n1584), .A(n978), .B(n977), .ZN(pc_out[13])
         );
  AOI22_X1 U1183 ( .A1(n233), .A2(\cache[0][1][DATA][12] ), .B1(n232), .B2(
        \cache[1][1][DATA][12] ), .ZN(n983) );
  AOI22_X1 U1184 ( .A1(n239), .A2(\cache[2][1][DATA][12] ), .B1(n37), .B2(
        \cache[3][1][DATA][12] ), .ZN(n982) );
  AOI22_X1 U1185 ( .A1(n243), .A2(\cache[4][1][DATA][12] ), .B1(n38), .B2(
        \cache[5][1][DATA][12] ), .ZN(n981) );
  AOI22_X1 U1186 ( .A1(n40), .A2(\cache[6][1][DATA][12] ), .B1(n39), .B2(
        \cache[7][1][DATA][12] ), .ZN(n980) );
  AND4_X1 U1187 ( .A1(n983), .A2(n982), .A3(n981), .A4(n980), .ZN(n1002) );
  AOI22_X1 U1188 ( .A1(n233), .A2(\cache[0][0][DATA][12] ), .B1(n232), .B2(
        \cache[1][0][DATA][12] ), .ZN(n987) );
  AOI22_X1 U1189 ( .A1(n240), .A2(\cache[2][0][DATA][12] ), .B1(n37), .B2(
        \cache[3][0][DATA][12] ), .ZN(n986) );
  AOI22_X1 U1190 ( .A1(n244), .A2(\cache[4][0][DATA][12] ), .B1(n38), .B2(
        \cache[5][0][DATA][12] ), .ZN(n985) );
  AOI22_X1 U1191 ( .A1(n40), .A2(\cache[6][0][DATA][12] ), .B1(n39), .B2(
        \cache[7][0][DATA][12] ), .ZN(n984) );
  NAND4_X1 U1192 ( .A1(n987), .A2(n986), .A3(n985), .A4(n984), .ZN(n994) );
  AOI22_X1 U1193 ( .A1(n235), .A2(\cache[0][2][DATA][12] ), .B1(n36), .B2(
        \cache[1][2][DATA][12] ), .ZN(n991) );
  AOI22_X1 U1194 ( .A1(n239), .A2(\cache[2][2][DATA][12] ), .B1(n37), .B2(
        \cache[3][2][DATA][12] ), .ZN(n990) );
  AOI22_X1 U1195 ( .A1(n243), .A2(\cache[4][2][DATA][12] ), .B1(n38), .B2(
        \cache[5][2][DATA][12] ), .ZN(n989) );
  AOI22_X1 U1196 ( .A1(n40), .A2(\cache[6][2][DATA][12] ), .B1(n39), .B2(
        \cache[7][2][DATA][12] ), .ZN(n988) );
  AND4_X1 U1197 ( .A1(n991), .A2(n990), .A3(n989), .A4(n988), .ZN(n992) );
  OAI22_X1 U1198 ( .A1(n992), .A2(n226), .B1(n275), .B2(n87), .ZN(n993) );
  AOI21_X1 U1199 ( .B1(n229), .B2(n994), .A(n993), .ZN(n1001) );
  AOI22_X1 U1200 ( .A1(n235), .A2(\cache[0][3][DATA][12] ), .B1(n36), .B2(
        \cache[1][3][DATA][12] ), .ZN(n998) );
  AOI22_X1 U1201 ( .A1(n55), .A2(\cache[2][3][DATA][12] ), .B1(n237), .B2(
        \cache[3][3][DATA][12] ), .ZN(n997) );
  AOI22_X1 U1202 ( .A1(n244), .A2(\cache[4][3][DATA][12] ), .B1(n241), .B2(
        \cache[5][3][DATA][12] ), .ZN(n996) );
  AOI22_X1 U1203 ( .A1(n40), .A2(\cache[6][3][DATA][12] ), .B1(n246), .B2(
        \cache[7][3][DATA][12] ), .ZN(n995) );
  NAND4_X1 U1204 ( .A1(n998), .A2(n997), .A3(n996), .A4(n995), .ZN(n999) );
  AOI22_X1 U1205 ( .A1(n248), .A2(n999), .B1(pc_in[14]), .B2(n93), .ZN(n1000)
         );
  OAI211_X1 U1206 ( .C1(n1002), .C2(n1584), .A(n1001), .B(n1000), .ZN(
        pc_out[14]) );
  AOI22_X1 U1207 ( .A1(n57), .A2(\cache[0][1][DATA][13] ), .B1(n36), .B2(
        \cache[1][1][DATA][13] ), .ZN(n1006) );
  AOI22_X1 U1208 ( .A1(n239), .A2(\cache[2][1][DATA][13] ), .B1(n37), .B2(
        \cache[3][1][DATA][13] ), .ZN(n1005) );
  AOI22_X1 U1209 ( .A1(n243), .A2(\cache[4][1][DATA][13] ), .B1(n38), .B2(
        \cache[5][1][DATA][13] ), .ZN(n1004) );
  AOI22_X1 U1210 ( .A1(n40), .A2(\cache[6][1][DATA][13] ), .B1(n246), .B2(
        \cache[7][1][DATA][13] ), .ZN(n1003) );
  AND4_X1 U1211 ( .A1(n1006), .A2(n1005), .A3(n1004), .A4(n1003), .ZN(n1025)
         );
  AOI22_X1 U1212 ( .A1(n236), .A2(\cache[0][0][DATA][13] ), .B1(n36), .B2(
        \cache[1][0][DATA][13] ), .ZN(n1010) );
  AOI22_X1 U1213 ( .A1(n239), .A2(\cache[2][0][DATA][13] ), .B1(n37), .B2(
        \cache[3][0][DATA][13] ), .ZN(n1009) );
  AOI22_X1 U1214 ( .A1(n243), .A2(\cache[4][0][DATA][13] ), .B1(n38), .B2(
        \cache[5][0][DATA][13] ), .ZN(n1008) );
  AOI22_X1 U1215 ( .A1(n40), .A2(\cache[6][0][DATA][13] ), .B1(n39), .B2(
        \cache[7][0][DATA][13] ), .ZN(n1007) );
  NAND4_X1 U1216 ( .A1(n1010), .A2(n1009), .A3(n1008), .A4(n1007), .ZN(n1017)
         );
  AOI22_X1 U1217 ( .A1(n236), .A2(\cache[0][2][DATA][13] ), .B1(n36), .B2(
        \cache[1][2][DATA][13] ), .ZN(n1014) );
  AOI22_X1 U1218 ( .A1(n240), .A2(\cache[2][2][DATA][13] ), .B1(n238), .B2(
        \cache[3][2][DATA][13] ), .ZN(n1013) );
  AOI22_X1 U1219 ( .A1(n244), .A2(\cache[4][2][DATA][13] ), .B1(n242), .B2(
        \cache[5][2][DATA][13] ), .ZN(n1012) );
  AOI22_X1 U1220 ( .A1(n40), .A2(\cache[6][2][DATA][13] ), .B1(n39), .B2(
        \cache[7][2][DATA][13] ), .ZN(n1011) );
  AND4_X1 U1221 ( .A1(n1014), .A2(n1013), .A3(n1012), .A4(n1011), .ZN(n1015)
         );
  OAI22_X1 U1222 ( .A1(n1015), .A2(n226), .B1(n276), .B2(n87), .ZN(n1016) );
  AOI21_X1 U1223 ( .B1(n230), .B2(n1017), .A(n1016), .ZN(n1024) );
  AOI22_X1 U1224 ( .A1(n57), .A2(\cache[0][3][DATA][13] ), .B1(n231), .B2(
        \cache[1][3][DATA][13] ), .ZN(n1021) );
  AOI22_X1 U1225 ( .A1(n240), .A2(\cache[2][3][DATA][13] ), .B1(n37), .B2(
        \cache[3][3][DATA][13] ), .ZN(n1020) );
  AOI22_X1 U1226 ( .A1(n244), .A2(\cache[4][3][DATA][13] ), .B1(n38), .B2(
        \cache[5][3][DATA][13] ), .ZN(n1019) );
  AOI22_X1 U1227 ( .A1(n40), .A2(\cache[6][3][DATA][13] ), .B1(n245), .B2(
        \cache[7][3][DATA][13] ), .ZN(n1018) );
  NAND4_X1 U1228 ( .A1(n1021), .A2(n1020), .A3(n1019), .A4(n1018), .ZN(n1022)
         );
  AOI22_X1 U1229 ( .A1(n248), .A2(n1022), .B1(pc_in[15]), .B2(n93), .ZN(n1023)
         );
  OAI211_X1 U1230 ( .C1(n1025), .C2(n1584), .A(n1024), .B(n1023), .ZN(
        pc_out[15]) );
  AOI22_X1 U1231 ( .A1(n57), .A2(\cache[0][1][DATA][14] ), .B1(n36), .B2(
        \cache[1][1][DATA][14] ), .ZN(n1029) );
  AOI22_X1 U1232 ( .A1(n240), .A2(\cache[2][1][DATA][14] ), .B1(n37), .B2(
        \cache[3][1][DATA][14] ), .ZN(n1028) );
  AOI22_X1 U1233 ( .A1(n244), .A2(\cache[4][1][DATA][14] ), .B1(n38), .B2(
        \cache[5][1][DATA][14] ), .ZN(n1027) );
  AOI22_X1 U1234 ( .A1(n40), .A2(\cache[6][1][DATA][14] ), .B1(n39), .B2(
        \cache[7][1][DATA][14] ), .ZN(n1026) );
  AND4_X1 U1235 ( .A1(n1029), .A2(n1028), .A3(n1027), .A4(n1026), .ZN(n1048)
         );
  AOI22_X1 U1236 ( .A1(n235), .A2(\cache[0][0][DATA][14] ), .B1(n36), .B2(
        \cache[1][0][DATA][14] ), .ZN(n1033) );
  AOI22_X1 U1237 ( .A1(n240), .A2(\cache[2][0][DATA][14] ), .B1(n238), .B2(
        \cache[3][0][DATA][14] ), .ZN(n1032) );
  AOI22_X1 U1238 ( .A1(n244), .A2(\cache[4][0][DATA][14] ), .B1(n38), .B2(
        \cache[5][0][DATA][14] ), .ZN(n1031) );
  AOI22_X1 U1239 ( .A1(n40), .A2(\cache[6][0][DATA][14] ), .B1(n39), .B2(
        \cache[7][0][DATA][14] ), .ZN(n1030) );
  NAND4_X1 U1240 ( .A1(n1033), .A2(n1032), .A3(n1031), .A4(n1030), .ZN(n1040)
         );
  AOI22_X1 U1241 ( .A1(n1569), .A2(\cache[0][2][DATA][14] ), .B1(n231), .B2(
        \cache[1][2][DATA][14] ), .ZN(n1037) );
  AOI22_X1 U1242 ( .A1(n240), .A2(\cache[2][2][DATA][14] ), .B1(n37), .B2(
        \cache[3][2][DATA][14] ), .ZN(n1036) );
  AOI22_X1 U1243 ( .A1(n244), .A2(\cache[4][2][DATA][14] ), .B1(n38), .B2(
        \cache[5][2][DATA][14] ), .ZN(n1035) );
  AOI22_X1 U1244 ( .A1(n40), .A2(\cache[6][2][DATA][14] ), .B1(n245), .B2(
        \cache[7][2][DATA][14] ), .ZN(n1034) );
  AND4_X1 U1245 ( .A1(n1037), .A2(n1036), .A3(n1035), .A4(n1034), .ZN(n1038)
         );
  OAI22_X1 U1246 ( .A1(n1038), .A2(n226), .B1(n277), .B2(n87), .ZN(n1039) );
  AOI21_X1 U1247 ( .B1(n26), .B2(n1040), .A(n1039), .ZN(n1047) );
  AOI22_X1 U1248 ( .A1(n57), .A2(\cache[0][3][DATA][14] ), .B1(n231), .B2(
        \cache[1][3][DATA][14] ), .ZN(n1044) );
  AOI22_X1 U1249 ( .A1(n240), .A2(\cache[2][3][DATA][14] ), .B1(n238), .B2(
        \cache[3][3][DATA][14] ), .ZN(n1043) );
  AOI22_X1 U1250 ( .A1(n244), .A2(\cache[4][3][DATA][14] ), .B1(n242), .B2(
        \cache[5][3][DATA][14] ), .ZN(n1042) );
  AOI22_X1 U1251 ( .A1(n40), .A2(\cache[6][3][DATA][14] ), .B1(n245), .B2(
        \cache[7][3][DATA][14] ), .ZN(n1041) );
  NAND4_X1 U1252 ( .A1(n1044), .A2(n1043), .A3(n1042), .A4(n1041), .ZN(n1045)
         );
  AOI22_X1 U1253 ( .A1(n96), .A2(n1045), .B1(pc_in[16]), .B2(n93), .ZN(n1046)
         );
  OAI211_X1 U1254 ( .C1(n1048), .C2(n1584), .A(n1047), .B(n1046), .ZN(
        pc_out[16]) );
  AOI22_X1 U1255 ( .A1(n233), .A2(\cache[0][1][DATA][15] ), .B1(n36), .B2(
        \cache[1][1][DATA][15] ), .ZN(n1052) );
  AOI22_X1 U1256 ( .A1(n240), .A2(\cache[2][1][DATA][15] ), .B1(n1570), .B2(
        \cache[3][1][DATA][15] ), .ZN(n1051) );
  AOI22_X1 U1257 ( .A1(n244), .A2(\cache[4][1][DATA][15] ), .B1(n1572), .B2(
        \cache[5][1][DATA][15] ), .ZN(n1050) );
  AOI22_X1 U1258 ( .A1(n40), .A2(\cache[6][1][DATA][15] ), .B1(n39), .B2(
        \cache[7][1][DATA][15] ), .ZN(n1049) );
  AND4_X1 U1259 ( .A1(n1052), .A2(n1051), .A3(n1050), .A4(n1049), .ZN(n1071)
         );
  AOI22_X1 U1260 ( .A1(n57), .A2(\cache[0][0][DATA][15] ), .B1(n36), .B2(
        \cache[1][0][DATA][15] ), .ZN(n1056) );
  AOI22_X1 U1261 ( .A1(n240), .A2(\cache[2][0][DATA][15] ), .B1(n238), .B2(
        \cache[3][0][DATA][15] ), .ZN(n1055) );
  AOI22_X1 U1262 ( .A1(n244), .A2(\cache[4][0][DATA][15] ), .B1(n38), .B2(
        \cache[5][0][DATA][15] ), .ZN(n1054) );
  AOI22_X1 U1263 ( .A1(n40), .A2(\cache[6][0][DATA][15] ), .B1(n39), .B2(
        \cache[7][0][DATA][15] ), .ZN(n1053) );
  NAND4_X1 U1264 ( .A1(n1056), .A2(n1055), .A3(n1054), .A4(n1053), .ZN(n1063)
         );
  AOI22_X1 U1265 ( .A1(n1569), .A2(\cache[0][2][DATA][15] ), .B1(n231), .B2(
        \cache[1][2][DATA][15] ), .ZN(n1060) );
  AOI22_X1 U1266 ( .A1(n240), .A2(\cache[2][2][DATA][15] ), .B1(n238), .B2(
        \cache[3][2][DATA][15] ), .ZN(n1059) );
  AOI22_X1 U1267 ( .A1(n244), .A2(\cache[4][2][DATA][15] ), .B1(n242), .B2(
        \cache[5][2][DATA][15] ), .ZN(n1058) );
  AOI22_X1 U1268 ( .A1(n40), .A2(\cache[6][2][DATA][15] ), .B1(n245), .B2(
        \cache[7][2][DATA][15] ), .ZN(n1057) );
  AND4_X1 U1269 ( .A1(n1060), .A2(n1059), .A3(n1058), .A4(n1057), .ZN(n1061)
         );
  OAI22_X1 U1270 ( .A1(n1061), .A2(n226), .B1(n278), .B2(n87), .ZN(n1062) );
  AOI21_X1 U1271 ( .B1(n229), .B2(n1063), .A(n1062), .ZN(n1070) );
  AOI22_X1 U1272 ( .A1(n233), .A2(\cache[0][3][DATA][15] ), .B1(n231), .B2(
        \cache[1][3][DATA][15] ), .ZN(n1067) );
  AOI22_X1 U1273 ( .A1(n240), .A2(\cache[2][3][DATA][15] ), .B1(n37), .B2(
        \cache[3][3][DATA][15] ), .ZN(n1066) );
  AOI22_X1 U1274 ( .A1(n244), .A2(\cache[4][3][DATA][15] ), .B1(n38), .B2(
        \cache[5][3][DATA][15] ), .ZN(n1065) );
  AOI22_X1 U1275 ( .A1(n40), .A2(\cache[6][3][DATA][15] ), .B1(n245), .B2(
        \cache[7][3][DATA][15] ), .ZN(n1064) );
  NAND4_X1 U1276 ( .A1(n1067), .A2(n1066), .A3(n1065), .A4(n1064), .ZN(n1068)
         );
  AOI22_X1 U1277 ( .A1(n248), .A2(n1068), .B1(pc_in[17]), .B2(n93), .ZN(n1069)
         );
  OAI211_X1 U1278 ( .C1(n1071), .C2(n1584), .A(n1070), .B(n1069), .ZN(
        pc_out[17]) );
  AOI22_X1 U1279 ( .A1(n57), .A2(\cache[0][1][DATA][16] ), .B1(n36), .B2(
        \cache[1][1][DATA][16] ), .ZN(n1075) );
  AOI22_X1 U1280 ( .A1(n240), .A2(\cache[2][1][DATA][16] ), .B1(n1570), .B2(
        \cache[3][1][DATA][16] ), .ZN(n1074) );
  AOI22_X1 U1281 ( .A1(n244), .A2(\cache[4][1][DATA][16] ), .B1(n1572), .B2(
        \cache[5][1][DATA][16] ), .ZN(n1073) );
  AOI22_X1 U1282 ( .A1(n40), .A2(\cache[6][1][DATA][16] ), .B1(n39), .B2(
        \cache[7][1][DATA][16] ), .ZN(n1072) );
  AND4_X1 U1283 ( .A1(n1075), .A2(n1074), .A3(n1073), .A4(n1072), .ZN(n1094)
         );
  AOI22_X1 U1284 ( .A1(n233), .A2(\cache[0][0][DATA][16] ), .B1(n36), .B2(
        \cache[1][0][DATA][16] ), .ZN(n1079) );
  AOI22_X1 U1285 ( .A1(n239), .A2(\cache[2][0][DATA][16] ), .B1(n37), .B2(
        \cache[3][0][DATA][16] ), .ZN(n1078) );
  AOI22_X1 U1286 ( .A1(n243), .A2(\cache[4][0][DATA][16] ), .B1(n242), .B2(
        \cache[5][0][DATA][16] ), .ZN(n1077) );
  AOI22_X1 U1287 ( .A1(n40), .A2(\cache[6][0][DATA][16] ), .B1(n39), .B2(
        \cache[7][0][DATA][16] ), .ZN(n1076) );
  NAND4_X1 U1288 ( .A1(n1079), .A2(n1078), .A3(n1077), .A4(n1076), .ZN(n1086)
         );
  AOI22_X1 U1289 ( .A1(n236), .A2(\cache[0][2][DATA][16] ), .B1(n232), .B2(
        \cache[1][2][DATA][16] ), .ZN(n1083) );
  AOI22_X1 U1290 ( .A1(n239), .A2(\cache[2][2][DATA][16] ), .B1(n237), .B2(
        \cache[3][2][DATA][16] ), .ZN(n1082) );
  AOI22_X1 U1291 ( .A1(n243), .A2(\cache[4][2][DATA][16] ), .B1(n241), .B2(
        \cache[5][2][DATA][16] ), .ZN(n1081) );
  AOI22_X1 U1292 ( .A1(n40), .A2(\cache[6][2][DATA][16] ), .B1(n39), .B2(
        \cache[7][2][DATA][16] ), .ZN(n1080) );
  AND4_X1 U1293 ( .A1(n1083), .A2(n1082), .A3(n1081), .A4(n1080), .ZN(n1084)
         );
  OAI22_X1 U1294 ( .A1(n1084), .A2(n226), .B1(n280), .B2(n88), .ZN(n1085) );
  AOI21_X1 U1295 ( .B1(n229), .B2(n1086), .A(n1085), .ZN(n1093) );
  AOI22_X1 U1296 ( .A1(n236), .A2(\cache[0][3][DATA][16] ), .B1(n232), .B2(
        \cache[1][3][DATA][16] ), .ZN(n1090) );
  AOI22_X1 U1297 ( .A1(n239), .A2(\cache[2][3][DATA][16] ), .B1(n237), .B2(
        \cache[3][3][DATA][16] ), .ZN(n1089) );
  AOI22_X1 U1298 ( .A1(n243), .A2(\cache[4][3][DATA][16] ), .B1(n241), .B2(
        \cache[5][3][DATA][16] ), .ZN(n1088) );
  AOI22_X1 U1299 ( .A1(n40), .A2(\cache[6][3][DATA][16] ), .B1(n246), .B2(
        \cache[7][3][DATA][16] ), .ZN(n1087) );
  NAND4_X1 U1300 ( .A1(n1090), .A2(n1089), .A3(n1088), .A4(n1087), .ZN(n1091)
         );
  AOI22_X1 U1301 ( .A1(n248), .A2(n1091), .B1(pc_in[18]), .B2(n93), .ZN(n1092)
         );
  OAI211_X1 U1302 ( .C1(n1094), .C2(n1584), .A(n1093), .B(n1092), .ZN(
        pc_out[18]) );
  AOI22_X1 U1303 ( .A1(n236), .A2(\cache[0][1][DATA][17] ), .B1(n232), .B2(
        \cache[1][1][DATA][17] ), .ZN(n1098) );
  AOI22_X1 U1304 ( .A1(n239), .A2(\cache[2][1][DATA][17] ), .B1(n37), .B2(
        \cache[3][1][DATA][17] ), .ZN(n1097) );
  AOI22_X1 U1305 ( .A1(n243), .A2(\cache[4][1][DATA][17] ), .B1(n38), .B2(
        \cache[5][1][DATA][17] ), .ZN(n1096) );
  AOI22_X1 U1306 ( .A1(n40), .A2(\cache[6][1][DATA][17] ), .B1(n246), .B2(
        \cache[7][1][DATA][17] ), .ZN(n1095) );
  AND4_X1 U1307 ( .A1(n1098), .A2(n1097), .A3(n1096), .A4(n1095), .ZN(n1117)
         );
  AOI22_X1 U1308 ( .A1(n236), .A2(\cache[0][0][DATA][17] ), .B1(n36), .B2(
        \cache[1][0][DATA][17] ), .ZN(n1102) );
  AOI22_X1 U1309 ( .A1(n239), .A2(\cache[2][0][DATA][17] ), .B1(n37), .B2(
        \cache[3][0][DATA][17] ), .ZN(n1101) );
  AOI22_X1 U1310 ( .A1(n243), .A2(\cache[4][0][DATA][17] ), .B1(n38), .B2(
        \cache[5][0][DATA][17] ), .ZN(n1100) );
  AOI22_X1 U1311 ( .A1(n40), .A2(\cache[6][0][DATA][17] ), .B1(n246), .B2(
        \cache[7][0][DATA][17] ), .ZN(n1099) );
  NAND4_X1 U1312 ( .A1(n1102), .A2(n1101), .A3(n1100), .A4(n1099), .ZN(n1109)
         );
  AOI22_X1 U1313 ( .A1(n236), .A2(\cache[0][2][DATA][17] ), .B1(n36), .B2(
        \cache[1][2][DATA][17] ), .ZN(n1106) );
  AOI22_X1 U1314 ( .A1(n239), .A2(\cache[2][2][DATA][17] ), .B1(n237), .B2(
        \cache[3][2][DATA][17] ), .ZN(n1105) );
  AOI22_X1 U1315 ( .A1(n243), .A2(\cache[4][2][DATA][17] ), .B1(n241), .B2(
        \cache[5][2][DATA][17] ), .ZN(n1104) );
  AOI22_X1 U1316 ( .A1(n40), .A2(\cache[6][2][DATA][17] ), .B1(n246), .B2(
        \cache[7][2][DATA][17] ), .ZN(n1103) );
  AND4_X1 U1317 ( .A1(n1106), .A2(n1105), .A3(n1104), .A4(n1103), .ZN(n1107)
         );
  OAI22_X1 U1318 ( .A1(n1107), .A2(n226), .B1(n281), .B2(n88), .ZN(n1108) );
  AOI21_X1 U1319 ( .B1(n230), .B2(n1109), .A(n1108), .ZN(n1116) );
  AOI22_X1 U1320 ( .A1(n236), .A2(\cache[0][3][DATA][17] ), .B1(n36), .B2(
        \cache[1][3][DATA][17] ), .ZN(n1113) );
  AOI22_X1 U1321 ( .A1(n239), .A2(\cache[2][3][DATA][17] ), .B1(n37), .B2(
        \cache[3][3][DATA][17] ), .ZN(n1112) );
  AOI22_X1 U1322 ( .A1(n243), .A2(\cache[4][3][DATA][17] ), .B1(n38), .B2(
        \cache[5][3][DATA][17] ), .ZN(n1111) );
  AOI22_X1 U1323 ( .A1(n40), .A2(\cache[6][3][DATA][17] ), .B1(n39), .B2(
        \cache[7][3][DATA][17] ), .ZN(n1110) );
  NAND4_X1 U1324 ( .A1(n1113), .A2(n1112), .A3(n1111), .A4(n1110), .ZN(n1114)
         );
  AOI22_X1 U1325 ( .A1(n248), .A2(n1114), .B1(pc_in[19]), .B2(n93), .ZN(n1115)
         );
  OAI211_X1 U1326 ( .C1(n1117), .C2(n1584), .A(n1116), .B(n1115), .ZN(
        pc_out[19]) );
  NAND2_X1 U1327 ( .A1(n1118), .A2(pc_in[1]), .ZN(n1119) );
  OAI21_X1 U1328 ( .B1(n1120), .B2(n88), .A(n1119), .ZN(pc_out[1]) );
  INV_X1 U1329 ( .A(pc_out[1]), .ZN(n585) );
  AOI22_X1 U1330 ( .A1(n236), .A2(\cache[0][1][DATA][18] ), .B1(n36), .B2(
        \cache[1][1][DATA][18] ), .ZN(n1124) );
  AOI22_X1 U1331 ( .A1(n239), .A2(\cache[2][1][DATA][18] ), .B1(n37), .B2(
        \cache[3][1][DATA][18] ), .ZN(n1123) );
  AOI22_X1 U1332 ( .A1(n243), .A2(\cache[4][1][DATA][18] ), .B1(n38), .B2(
        \cache[5][1][DATA][18] ), .ZN(n1122) );
  AOI22_X1 U1333 ( .A1(n40), .A2(\cache[6][1][DATA][18] ), .B1(n246), .B2(
        \cache[7][1][DATA][18] ), .ZN(n1121) );
  AND4_X1 U1334 ( .A1(n1124), .A2(n1123), .A3(n1122), .A4(n1121), .ZN(n1143)
         );
  AOI22_X1 U1335 ( .A1(n236), .A2(\cache[0][0][DATA][18] ), .B1(n232), .B2(
        \cache[1][0][DATA][18] ), .ZN(n1128) );
  AOI22_X1 U1336 ( .A1(n239), .A2(\cache[2][0][DATA][18] ), .B1(n37), .B2(
        \cache[3][0][DATA][18] ), .ZN(n1127) );
  AOI22_X1 U1337 ( .A1(n243), .A2(\cache[4][0][DATA][18] ), .B1(n38), .B2(
        \cache[5][0][DATA][18] ), .ZN(n1126) );
  AOI22_X1 U1338 ( .A1(n40), .A2(\cache[6][0][DATA][18] ), .B1(n39), .B2(
        \cache[7][0][DATA][18] ), .ZN(n1125) );
  NAND4_X1 U1339 ( .A1(n1128), .A2(n1127), .A3(n1126), .A4(n1125), .ZN(n1135)
         );
  AOI22_X1 U1340 ( .A1(n236), .A2(\cache[0][2][DATA][18] ), .B1(n232), .B2(
        \cache[1][2][DATA][18] ), .ZN(n1132) );
  AOI22_X1 U1341 ( .A1(n239), .A2(\cache[2][2][DATA][18] ), .B1(n237), .B2(
        \cache[3][2][DATA][18] ), .ZN(n1131) );
  AOI22_X1 U1342 ( .A1(n243), .A2(\cache[4][2][DATA][18] ), .B1(n241), .B2(
        \cache[5][2][DATA][18] ), .ZN(n1130) );
  AOI22_X1 U1343 ( .A1(n40), .A2(\cache[6][2][DATA][18] ), .B1(n39), .B2(
        \cache[7][2][DATA][18] ), .ZN(n1129) );
  AND4_X1 U1344 ( .A1(n1132), .A2(n1131), .A3(n1130), .A4(n1129), .ZN(n1133)
         );
  OAI22_X1 U1345 ( .A1(n1133), .A2(n226), .B1(n282), .B2(n88), .ZN(n1134) );
  AOI21_X1 U1346 ( .B1(n229), .B2(n1135), .A(n1134), .ZN(n1142) );
  AOI22_X1 U1347 ( .A1(n236), .A2(\cache[0][3][DATA][18] ), .B1(n232), .B2(
        \cache[1][3][DATA][18] ), .ZN(n1139) );
  AOI22_X1 U1348 ( .A1(n239), .A2(\cache[2][3][DATA][18] ), .B1(n237), .B2(
        \cache[3][3][DATA][18] ), .ZN(n1138) );
  AOI22_X1 U1349 ( .A1(n243), .A2(\cache[4][3][DATA][18] ), .B1(n241), .B2(
        \cache[5][3][DATA][18] ), .ZN(n1137) );
  AOI22_X1 U1350 ( .A1(n40), .A2(\cache[6][3][DATA][18] ), .B1(n39), .B2(
        \cache[7][3][DATA][18] ), .ZN(n1136) );
  NAND4_X1 U1351 ( .A1(n1139), .A2(n1138), .A3(n1137), .A4(n1136), .ZN(n1140)
         );
  AOI22_X1 U1352 ( .A1(n248), .A2(n1140), .B1(pc_in[20]), .B2(n93), .ZN(n1141)
         );
  OAI211_X1 U1353 ( .C1(n1143), .C2(n1584), .A(n1142), .B(n1141), .ZN(
        pc_out[20]) );
  AOI22_X1 U1354 ( .A1(n235), .A2(\cache[0][1][DATA][19] ), .B1(n36), .B2(
        \cache[1][1][DATA][19] ), .ZN(n1147) );
  AOI22_X1 U1355 ( .A1(n239), .A2(\cache[2][1][DATA][19] ), .B1(n1570), .B2(
        \cache[3][1][DATA][19] ), .ZN(n1146) );
  AOI22_X1 U1356 ( .A1(n243), .A2(\cache[4][1][DATA][19] ), .B1(n38), .B2(
        \cache[5][1][DATA][19] ), .ZN(n1145) );
  AOI22_X1 U1357 ( .A1(n40), .A2(\cache[6][1][DATA][19] ), .B1(n39), .B2(
        \cache[7][1][DATA][19] ), .ZN(n1144) );
  AND4_X1 U1358 ( .A1(n1147), .A2(n1146), .A3(n1145), .A4(n1144), .ZN(n1166)
         );
  AOI22_X1 U1359 ( .A1(n235), .A2(\cache[0][0][DATA][19] ), .B1(n36), .B2(
        \cache[1][0][DATA][19] ), .ZN(n1151) );
  AOI22_X1 U1360 ( .A1(n239), .A2(\cache[2][0][DATA][19] ), .B1(n37), .B2(
        \cache[3][0][DATA][19] ), .ZN(n1150) );
  AOI22_X1 U1361 ( .A1(n243), .A2(\cache[4][0][DATA][19] ), .B1(n242), .B2(
        \cache[5][0][DATA][19] ), .ZN(n1149) );
  AOI22_X1 U1362 ( .A1(n40), .A2(\cache[6][0][DATA][19] ), .B1(n39), .B2(
        \cache[7][0][DATA][19] ), .ZN(n1148) );
  NAND4_X1 U1363 ( .A1(n1151), .A2(n1150), .A3(n1149), .A4(n1148), .ZN(n1158)
         );
  AOI22_X1 U1364 ( .A1(n235), .A2(\cache[0][2][DATA][19] ), .B1(n36), .B2(
        \cache[1][2][DATA][19] ), .ZN(n1155) );
  AOI22_X1 U1365 ( .A1(n239), .A2(\cache[2][2][DATA][19] ), .B1(n37), .B2(
        \cache[3][2][DATA][19] ), .ZN(n1154) );
  AOI22_X1 U1366 ( .A1(n243), .A2(\cache[4][2][DATA][19] ), .B1(n38), .B2(
        \cache[5][2][DATA][19] ), .ZN(n1153) );
  AOI22_X1 U1367 ( .A1(n40), .A2(\cache[6][2][DATA][19] ), .B1(n39), .B2(
        \cache[7][2][DATA][19] ), .ZN(n1152) );
  AND4_X1 U1368 ( .A1(n1155), .A2(n1154), .A3(n1153), .A4(n1152), .ZN(n1156)
         );
  OAI22_X1 U1369 ( .A1(n1156), .A2(n226), .B1(n283), .B2(n88), .ZN(n1157) );
  AOI21_X1 U1370 ( .B1(n230), .B2(n1158), .A(n1157), .ZN(n1165) );
  AOI22_X1 U1371 ( .A1(n235), .A2(\cache[0][3][DATA][19] ), .B1(n231), .B2(
        \cache[1][3][DATA][19] ), .ZN(n1162) );
  AOI22_X1 U1372 ( .A1(n239), .A2(\cache[2][3][DATA][19] ), .B1(n37), .B2(
        \cache[3][3][DATA][19] ), .ZN(n1161) );
  AOI22_X1 U1373 ( .A1(n243), .A2(\cache[4][3][DATA][19] ), .B1(n38), .B2(
        \cache[5][3][DATA][19] ), .ZN(n1160) );
  AOI22_X1 U1374 ( .A1(n40), .A2(\cache[6][3][DATA][19] ), .B1(n245), .B2(
        \cache[7][3][DATA][19] ), .ZN(n1159) );
  NAND4_X1 U1375 ( .A1(n1162), .A2(n1161), .A3(n1160), .A4(n1159), .ZN(n1163)
         );
  AOI22_X1 U1376 ( .A1(n248), .A2(n1163), .B1(pc_in[21]), .B2(n91), .ZN(n1164)
         );
  OAI211_X1 U1377 ( .C1(n1166), .C2(n1584), .A(n1165), .B(n1164), .ZN(
        pc_out[21]) );
  AOI22_X1 U1378 ( .A1(n235), .A2(\cache[0][1][DATA][20] ), .B1(n36), .B2(
        \cache[1][1][DATA][20] ), .ZN(n1170) );
  AOI22_X1 U1379 ( .A1(n239), .A2(\cache[2][1][DATA][20] ), .B1(n37), .B2(
        \cache[3][1][DATA][20] ), .ZN(n1169) );
  AOI22_X1 U1380 ( .A1(n243), .A2(\cache[4][1][DATA][20] ), .B1(n1572), .B2(
        \cache[5][1][DATA][20] ), .ZN(n1168) );
  AOI22_X1 U1381 ( .A1(n40), .A2(\cache[6][1][DATA][20] ), .B1(n39), .B2(
        \cache[7][1][DATA][20] ), .ZN(n1167) );
  AND4_X1 U1382 ( .A1(n1170), .A2(n1169), .A3(n1168), .A4(n1167), .ZN(n1189)
         );
  AOI22_X1 U1383 ( .A1(n235), .A2(\cache[0][0][DATA][20] ), .B1(n36), .B2(
        \cache[1][0][DATA][20] ), .ZN(n1174) );
  AOI22_X1 U1384 ( .A1(n239), .A2(\cache[2][0][DATA][20] ), .B1(n37), .B2(
        \cache[3][0][DATA][20] ), .ZN(n1173) );
  AOI22_X1 U1385 ( .A1(n243), .A2(\cache[4][0][DATA][20] ), .B1(n38), .B2(
        \cache[5][0][DATA][20] ), .ZN(n1172) );
  AOI22_X1 U1386 ( .A1(n40), .A2(\cache[6][0][DATA][20] ), .B1(n39), .B2(
        \cache[7][0][DATA][20] ), .ZN(n1171) );
  NAND4_X1 U1387 ( .A1(n1174), .A2(n1173), .A3(n1172), .A4(n1171), .ZN(n1181)
         );
  AOI22_X1 U1388 ( .A1(n235), .A2(\cache[0][2][DATA][20] ), .B1(n36), .B2(
        \cache[1][2][DATA][20] ), .ZN(n1178) );
  AOI22_X1 U1389 ( .A1(n239), .A2(\cache[2][2][DATA][20] ), .B1(n238), .B2(
        \cache[3][2][DATA][20] ), .ZN(n1177) );
  AOI22_X1 U1390 ( .A1(n243), .A2(\cache[4][2][DATA][20] ), .B1(n242), .B2(
        \cache[5][2][DATA][20] ), .ZN(n1176) );
  AOI22_X1 U1391 ( .A1(n40), .A2(\cache[6][2][DATA][20] ), .B1(n39), .B2(
        \cache[7][2][DATA][20] ), .ZN(n1175) );
  AND4_X1 U1392 ( .A1(n1178), .A2(n1177), .A3(n1176), .A4(n1175), .ZN(n1179)
         );
  OAI22_X1 U1393 ( .A1(n1179), .A2(n226), .B1(n284), .B2(n88), .ZN(n1180) );
  AOI21_X1 U1394 ( .B1(n229), .B2(n1181), .A(n1180), .ZN(n1188) );
  AOI22_X1 U1395 ( .A1(n235), .A2(\cache[0][3][DATA][20] ), .B1(n231), .B2(
        \cache[1][3][DATA][20] ), .ZN(n1185) );
  AOI22_X1 U1396 ( .A1(n239), .A2(\cache[2][3][DATA][20] ), .B1(n37), .B2(
        \cache[3][3][DATA][20] ), .ZN(n1184) );
  AOI22_X1 U1397 ( .A1(n243), .A2(\cache[4][3][DATA][20] ), .B1(n38), .B2(
        \cache[5][3][DATA][20] ), .ZN(n1183) );
  AOI22_X1 U1398 ( .A1(n40), .A2(\cache[6][3][DATA][20] ), .B1(n245), .B2(
        \cache[7][3][DATA][20] ), .ZN(n1182) );
  NAND4_X1 U1399 ( .A1(n1185), .A2(n1184), .A3(n1183), .A4(n1182), .ZN(n1186)
         );
  AOI22_X1 U1400 ( .A1(n248), .A2(n1186), .B1(pc_in[22]), .B2(n91), .ZN(n1187)
         );
  OAI211_X1 U1401 ( .C1(n1189), .C2(n1584), .A(n1188), .B(n1187), .ZN(
        pc_out[22]) );
  AOI22_X1 U1402 ( .A1(n235), .A2(\cache[0][1][DATA][21] ), .B1(n36), .B2(
        \cache[1][1][DATA][21] ), .ZN(n1193) );
  AOI22_X1 U1403 ( .A1(n239), .A2(\cache[2][1][DATA][21] ), .B1(n238), .B2(
        \cache[3][1][DATA][21] ), .ZN(n1192) );
  AOI22_X1 U1404 ( .A1(n243), .A2(\cache[4][1][DATA][21] ), .B1(n242), .B2(
        \cache[5][1][DATA][21] ), .ZN(n1191) );
  AOI22_X1 U1405 ( .A1(n40), .A2(\cache[6][1][DATA][21] ), .B1(n39), .B2(
        \cache[7][1][DATA][21] ), .ZN(n1190) );
  AND4_X1 U1406 ( .A1(n1193), .A2(n1192), .A3(n1191), .A4(n1190), .ZN(n1212)
         );
  AOI22_X1 U1407 ( .A1(n235), .A2(\cache[0][0][DATA][21] ), .B1(n36), .B2(
        \cache[1][0][DATA][21] ), .ZN(n1197) );
  AOI22_X1 U1408 ( .A1(n239), .A2(\cache[2][0][DATA][21] ), .B1(n238), .B2(
        \cache[3][0][DATA][21] ), .ZN(n1196) );
  AOI22_X1 U1409 ( .A1(n243), .A2(\cache[4][0][DATA][21] ), .B1(n242), .B2(
        \cache[5][0][DATA][21] ), .ZN(n1195) );
  AOI22_X1 U1410 ( .A1(n40), .A2(\cache[6][0][DATA][21] ), .B1(n39), .B2(
        \cache[7][0][DATA][21] ), .ZN(n1194) );
  NAND4_X1 U1411 ( .A1(n1197), .A2(n1196), .A3(n1195), .A4(n1194), .ZN(n1204)
         );
  AOI22_X1 U1412 ( .A1(n235), .A2(\cache[0][2][DATA][21] ), .B1(n36), .B2(
        \cache[1][2][DATA][21] ), .ZN(n1201) );
  AOI22_X1 U1413 ( .A1(n55), .A2(\cache[2][2][DATA][21] ), .B1(n37), .B2(
        \cache[3][2][DATA][21] ), .ZN(n1200) );
  AOI22_X1 U1414 ( .A1(n56), .A2(\cache[4][2][DATA][21] ), .B1(n38), .B2(
        \cache[5][2][DATA][21] ), .ZN(n1199) );
  AOI22_X1 U1415 ( .A1(n40), .A2(\cache[6][2][DATA][21] ), .B1(n39), .B2(
        \cache[7][2][DATA][21] ), .ZN(n1198) );
  AND4_X1 U1416 ( .A1(n1201), .A2(n1200), .A3(n1199), .A4(n1198), .ZN(n1202)
         );
  OAI22_X1 U1417 ( .A1(n1202), .A2(n226), .B1(n285), .B2(n88), .ZN(n1203) );
  AOI21_X1 U1418 ( .B1(n230), .B2(n1204), .A(n1203), .ZN(n1211) );
  AOI22_X1 U1419 ( .A1(n234), .A2(\cache[0][3][DATA][21] ), .B1(n36), .B2(
        \cache[1][3][DATA][21] ), .ZN(n1208) );
  AOI22_X1 U1420 ( .A1(n55), .A2(\cache[2][3][DATA][21] ), .B1(n37), .B2(
        \cache[3][3][DATA][21] ), .ZN(n1207) );
  AOI22_X1 U1421 ( .A1(n56), .A2(\cache[4][3][DATA][21] ), .B1(n38), .B2(
        \cache[5][3][DATA][21] ), .ZN(n1206) );
  AOI22_X1 U1422 ( .A1(n40), .A2(\cache[6][3][DATA][21] ), .B1(n39), .B2(
        \cache[7][3][DATA][21] ), .ZN(n1205) );
  NAND4_X1 U1423 ( .A1(n1208), .A2(n1207), .A3(n1206), .A4(n1205), .ZN(n1209)
         );
  AOI22_X1 U1424 ( .A1(n96), .A2(n1209), .B1(pc_in[23]), .B2(n93), .ZN(n1210)
         );
  OAI211_X1 U1425 ( .C1(n1212), .C2(n1584), .A(n1211), .B(n1210), .ZN(
        pc_out[23]) );
  AOI22_X1 U1426 ( .A1(n234), .A2(\cache[0][1][DATA][22] ), .B1(n36), .B2(
        \cache[1][1][DATA][22] ), .ZN(n1216) );
  AOI22_X1 U1427 ( .A1(n55), .A2(\cache[2][1][DATA][22] ), .B1(n37), .B2(
        \cache[3][1][DATA][22] ), .ZN(n1215) );
  AOI22_X1 U1428 ( .A1(n56), .A2(\cache[4][1][DATA][22] ), .B1(n38), .B2(
        \cache[5][1][DATA][22] ), .ZN(n1214) );
  AOI22_X1 U1429 ( .A1(n40), .A2(\cache[6][1][DATA][22] ), .B1(n39), .B2(
        \cache[7][1][DATA][22] ), .ZN(n1213) );
  AND4_X1 U1430 ( .A1(n1216), .A2(n1215), .A3(n1214), .A4(n1213), .ZN(n1235)
         );
  AOI22_X1 U1431 ( .A1(n234), .A2(\cache[0][0][DATA][22] ), .B1(n231), .B2(
        \cache[1][0][DATA][22] ), .ZN(n1220) );
  AOI22_X1 U1432 ( .A1(n55), .A2(\cache[2][0][DATA][22] ), .B1(n237), .B2(
        \cache[3][0][DATA][22] ), .ZN(n1219) );
  AOI22_X1 U1433 ( .A1(n56), .A2(\cache[4][0][DATA][22] ), .B1(n241), .B2(
        \cache[5][0][DATA][22] ), .ZN(n1218) );
  AOI22_X1 U1434 ( .A1(n40), .A2(\cache[6][0][DATA][22] ), .B1(n245), .B2(
        \cache[7][0][DATA][22] ), .ZN(n1217) );
  NAND4_X1 U1435 ( .A1(n1220), .A2(n1219), .A3(n1218), .A4(n1217), .ZN(n1227)
         );
  AOI22_X1 U1436 ( .A1(n234), .A2(\cache[0][2][DATA][22] ), .B1(n231), .B2(
        \cache[1][2][DATA][22] ), .ZN(n1224) );
  AOI22_X1 U1437 ( .A1(n55), .A2(\cache[2][2][DATA][22] ), .B1(n237), .B2(
        \cache[3][2][DATA][22] ), .ZN(n1223) );
  AOI22_X1 U1438 ( .A1(n56), .A2(\cache[4][2][DATA][22] ), .B1(n241), .B2(
        \cache[5][2][DATA][22] ), .ZN(n1222) );
  AOI22_X1 U1439 ( .A1(n40), .A2(\cache[6][2][DATA][22] ), .B1(n245), .B2(
        \cache[7][2][DATA][22] ), .ZN(n1221) );
  AND4_X1 U1440 ( .A1(n1224), .A2(n1223), .A3(n1222), .A4(n1221), .ZN(n1225)
         );
  AOI22_X1 U1441 ( .A1(n234), .A2(\cache[0][3][DATA][22] ), .B1(n231), .B2(
        \cache[1][3][DATA][22] ), .ZN(n1231) );
  AOI22_X1 U1442 ( .A1(n55), .A2(\cache[2][3][DATA][22] ), .B1(n237), .B2(
        \cache[3][3][DATA][22] ), .ZN(n1230) );
  AOI22_X1 U1443 ( .A1(n56), .A2(\cache[4][3][DATA][22] ), .B1(n241), .B2(
        \cache[5][3][DATA][22] ), .ZN(n1229) );
  AOI22_X1 U1444 ( .A1(n40), .A2(\cache[6][3][DATA][22] ), .B1(n245), .B2(
        \cache[7][3][DATA][22] ), .ZN(n1228) );
  NAND4_X1 U1445 ( .A1(n1231), .A2(n1230), .A3(n1229), .A4(n1228), .ZN(n1232)
         );
  AOI22_X1 U1446 ( .A1(n249), .A2(n1232), .B1(pc_in[24]), .B2(n93), .ZN(n1233)
         );
  OAI211_X1 U1447 ( .C1(n1235), .C2(n1584), .A(n1233), .B(n1234), .ZN(
        pc_out[24]) );
  AOI22_X1 U1448 ( .A1(n234), .A2(\cache[0][1][DATA][23] ), .B1(n36), .B2(
        \cache[1][1][DATA][23] ), .ZN(n1239) );
  AOI22_X1 U1449 ( .A1(n55), .A2(\cache[2][1][DATA][23] ), .B1(n37), .B2(
        \cache[3][1][DATA][23] ), .ZN(n1238) );
  AOI22_X1 U1450 ( .A1(n56), .A2(\cache[4][1][DATA][23] ), .B1(n38), .B2(
        \cache[5][1][DATA][23] ), .ZN(n1237) );
  AOI22_X1 U1451 ( .A1(n40), .A2(\cache[6][1][DATA][23] ), .B1(n39), .B2(
        \cache[7][1][DATA][23] ), .ZN(n1236) );
  AND4_X1 U1452 ( .A1(n1239), .A2(n1238), .A3(n1237), .A4(n1236), .ZN(n1258)
         );
  AOI22_X1 U1453 ( .A1(n234), .A2(\cache[0][0][DATA][23] ), .B1(n36), .B2(
        \cache[1][0][DATA][23] ), .ZN(n1243) );
  AOI22_X1 U1454 ( .A1(n55), .A2(\cache[2][0][DATA][23] ), .B1(n237), .B2(
        \cache[3][0][DATA][23] ), .ZN(n1242) );
  AOI22_X1 U1455 ( .A1(n56), .A2(\cache[4][0][DATA][23] ), .B1(n241), .B2(
        \cache[5][0][DATA][23] ), .ZN(n1241) );
  AOI22_X1 U1456 ( .A1(n40), .A2(\cache[6][0][DATA][23] ), .B1(n245), .B2(
        \cache[7][0][DATA][23] ), .ZN(n1240) );
  NAND4_X1 U1457 ( .A1(n1243), .A2(n1242), .A3(n1241), .A4(n1240), .ZN(n1250)
         );
  AOI22_X1 U1458 ( .A1(n234), .A2(\cache[0][2][DATA][23] ), .B1(n231), .B2(
        \cache[1][2][DATA][23] ), .ZN(n1247) );
  AOI22_X1 U1459 ( .A1(n55), .A2(\cache[2][2][DATA][23] ), .B1(n237), .B2(
        \cache[3][2][DATA][23] ), .ZN(n1246) );
  AOI22_X1 U1460 ( .A1(n56), .A2(\cache[4][2][DATA][23] ), .B1(n241), .B2(
        \cache[5][2][DATA][23] ), .ZN(n1245) );
  AOI22_X1 U1461 ( .A1(n40), .A2(\cache[6][2][DATA][23] ), .B1(n245), .B2(
        \cache[7][2][DATA][23] ), .ZN(n1244) );
  AND4_X1 U1462 ( .A1(n1247), .A2(n1246), .A3(n1245), .A4(n1244), .ZN(n1248)
         );
  AOI22_X1 U1463 ( .A1(n234), .A2(\cache[0][3][DATA][23] ), .B1(n231), .B2(
        \cache[1][3][DATA][23] ), .ZN(n1254) );
  AOI22_X1 U1464 ( .A1(n55), .A2(\cache[2][3][DATA][23] ), .B1(n237), .B2(
        \cache[3][3][DATA][23] ), .ZN(n1253) );
  AOI22_X1 U1465 ( .A1(n56), .A2(\cache[4][3][DATA][23] ), .B1(n241), .B2(
        \cache[5][3][DATA][23] ), .ZN(n1252) );
  AOI22_X1 U1466 ( .A1(n40), .A2(\cache[6][3][DATA][23] ), .B1(n245), .B2(
        \cache[7][3][DATA][23] ), .ZN(n1251) );
  NAND4_X1 U1467 ( .A1(n1254), .A2(n1253), .A3(n1252), .A4(n1251), .ZN(n1255)
         );
  AOI22_X1 U1468 ( .A1(n96), .A2(n1255), .B1(pc_in[25]), .B2(n93), .ZN(n1256)
         );
  OAI211_X1 U1469 ( .C1(n1258), .C2(n1584), .A(n1257), .B(n1256), .ZN(
        pc_out[25]) );
  AOI22_X1 U1470 ( .A1(n234), .A2(\cache[0][1][DATA][24] ), .B1(n36), .B2(
        \cache[1][1][DATA][24] ), .ZN(n1262) );
  AOI22_X1 U1471 ( .A1(n55), .A2(\cache[2][1][DATA][24] ), .B1(n37), .B2(
        \cache[3][1][DATA][24] ), .ZN(n1261) );
  AOI22_X1 U1472 ( .A1(n56), .A2(\cache[4][1][DATA][24] ), .B1(n38), .B2(
        \cache[5][1][DATA][24] ), .ZN(n1260) );
  AOI22_X1 U1473 ( .A1(n40), .A2(\cache[6][1][DATA][24] ), .B1(n39), .B2(
        \cache[7][1][DATA][24] ), .ZN(n1259) );
  AND4_X1 U1474 ( .A1(n1262), .A2(n1261), .A3(n1260), .A4(n1259), .ZN(n1281)
         );
  AOI22_X1 U1475 ( .A1(n234), .A2(\cache[0][0][DATA][24] ), .B1(n36), .B2(
        \cache[1][0][DATA][24] ), .ZN(n1266) );
  AOI22_X1 U1476 ( .A1(n239), .A2(\cache[2][0][DATA][24] ), .B1(n37), .B2(
        \cache[3][0][DATA][24] ), .ZN(n1265) );
  AOI22_X1 U1477 ( .A1(n56), .A2(\cache[4][0][DATA][24] ), .B1(n38), .B2(
        \cache[5][0][DATA][24] ), .ZN(n1264) );
  AOI22_X1 U1478 ( .A1(n40), .A2(\cache[6][0][DATA][24] ), .B1(n39), .B2(
        \cache[7][0][DATA][24] ), .ZN(n1263) );
  NAND4_X1 U1479 ( .A1(n1266), .A2(n1265), .A3(n1264), .A4(n1263), .ZN(n1273)
         );
  AOI22_X1 U1480 ( .A1(n233), .A2(\cache[0][2][DATA][24] ), .B1(n231), .B2(
        \cache[1][2][DATA][24] ), .ZN(n1270) );
  AOI22_X1 U1481 ( .A1(n240), .A2(\cache[2][2][DATA][24] ), .B1(n37), .B2(
        \cache[3][2][DATA][24] ), .ZN(n1269) );
  AOI22_X1 U1482 ( .A1(n244), .A2(\cache[4][2][DATA][24] ), .B1(n38), .B2(
        \cache[5][2][DATA][24] ), .ZN(n1268) );
  AOI22_X1 U1483 ( .A1(n40), .A2(\cache[6][2][DATA][24] ), .B1(n39), .B2(
        \cache[7][2][DATA][24] ), .ZN(n1267) );
  AND4_X1 U1484 ( .A1(n1270), .A2(n1269), .A3(n1268), .A4(n1267), .ZN(n1271)
         );
  AOI21_X1 U1485 ( .B1(n230), .B2(n1273), .A(n1272), .ZN(n1280) );
  AOI22_X1 U1486 ( .A1(n233), .A2(\cache[0][3][DATA][24] ), .B1(n36), .B2(
        \cache[1][3][DATA][24] ), .ZN(n1277) );
  AOI22_X1 U1487 ( .A1(n240), .A2(\cache[2][3][DATA][24] ), .B1(n37), .B2(
        \cache[3][3][DATA][24] ), .ZN(n1276) );
  AOI22_X1 U1488 ( .A1(n244), .A2(\cache[4][3][DATA][24] ), .B1(n38), .B2(
        \cache[5][3][DATA][24] ), .ZN(n1275) );
  AOI22_X1 U1489 ( .A1(n40), .A2(\cache[6][3][DATA][24] ), .B1(n39), .B2(
        \cache[7][3][DATA][24] ), .ZN(n1274) );
  NAND4_X1 U1490 ( .A1(n1277), .A2(n1276), .A3(n1275), .A4(n1274), .ZN(n1278)
         );
  AOI22_X1 U1491 ( .A1(n249), .A2(n1278), .B1(pc_in[26]), .B2(n93), .ZN(n1279)
         );
  AOI22_X1 U1492 ( .A1(n233), .A2(\cache[0][1][DATA][25] ), .B1(n231), .B2(
        \cache[1][1][DATA][25] ), .ZN(n1285) );
  AOI22_X1 U1493 ( .A1(n239), .A2(\cache[2][1][DATA][25] ), .B1(n237), .B2(
        \cache[3][1][DATA][25] ), .ZN(n1284) );
  AOI22_X1 U1494 ( .A1(n56), .A2(\cache[4][1][DATA][25] ), .B1(n241), .B2(
        \cache[5][1][DATA][25] ), .ZN(n1283) );
  AOI22_X1 U1495 ( .A1(n40), .A2(\cache[6][1][DATA][25] ), .B1(n245), .B2(
        \cache[7][1][DATA][25] ), .ZN(n1282) );
  AND4_X1 U1496 ( .A1(n1285), .A2(n1284), .A3(n1283), .A4(n1282), .ZN(n1304)
         );
  AOI22_X1 U1497 ( .A1(n233), .A2(\cache[0][0][DATA][25] ), .B1(n36), .B2(
        \cache[1][0][DATA][25] ), .ZN(n1289) );
  AOI22_X1 U1498 ( .A1(n55), .A2(\cache[2][0][DATA][25] ), .B1(n37), .B2(
        \cache[3][0][DATA][25] ), .ZN(n1288) );
  AOI22_X1 U1499 ( .A1(n244), .A2(\cache[4][0][DATA][25] ), .B1(n38), .B2(
        \cache[5][0][DATA][25] ), .ZN(n1287) );
  AOI22_X1 U1500 ( .A1(n40), .A2(\cache[6][0][DATA][25] ), .B1(n39), .B2(
        \cache[7][0][DATA][25] ), .ZN(n1286) );
  NAND4_X1 U1501 ( .A1(n1289), .A2(n1288), .A3(n1287), .A4(n1286), .ZN(n1296)
         );
  AOI22_X1 U1502 ( .A1(n233), .A2(\cache[0][2][DATA][25] ), .B1(n36), .B2(
        \cache[1][2][DATA][25] ), .ZN(n1293) );
  AOI22_X1 U1503 ( .A1(n55), .A2(\cache[2][2][DATA][25] ), .B1(n37), .B2(
        \cache[3][2][DATA][25] ), .ZN(n1292) );
  AOI22_X1 U1504 ( .A1(n56), .A2(\cache[4][2][DATA][25] ), .B1(n38), .B2(
        \cache[5][2][DATA][25] ), .ZN(n1291) );
  AOI22_X1 U1505 ( .A1(n40), .A2(\cache[6][2][DATA][25] ), .B1(n39), .B2(
        \cache[7][2][DATA][25] ), .ZN(n1290) );
  AND4_X1 U1506 ( .A1(n1293), .A2(n1292), .A3(n1291), .A4(n1290), .ZN(n1294)
         );
  AOI22_X1 U1507 ( .A1(n233), .A2(\cache[0][3][DATA][25] ), .B1(n36), .B2(
        \cache[1][3][DATA][25] ), .ZN(n1300) );
  AOI22_X1 U1508 ( .A1(n240), .A2(\cache[2][3][DATA][25] ), .B1(n37), .B2(
        \cache[3][3][DATA][25] ), .ZN(n1299) );
  AOI22_X1 U1509 ( .A1(n244), .A2(\cache[4][3][DATA][25] ), .B1(n38), .B2(
        \cache[5][3][DATA][25] ), .ZN(n1298) );
  AOI22_X1 U1510 ( .A1(n40), .A2(\cache[6][3][DATA][25] ), .B1(n39), .B2(
        \cache[7][3][DATA][25] ), .ZN(n1297) );
  NAND4_X1 U1511 ( .A1(n1300), .A2(n1299), .A3(n1298), .A4(n1297), .ZN(n1301)
         );
  AOI22_X1 U1512 ( .A1(n96), .A2(n1301), .B1(pc_in[27]), .B2(n91), .ZN(n1302)
         );
  OAI211_X1 U1513 ( .C1(n1304), .C2(n1584), .A(n1303), .B(n1302), .ZN(
        pc_out[27]) );
  AOI22_X1 U1514 ( .A1(n233), .A2(\cache[0][1][DATA][26] ), .B1(n231), .B2(
        \cache[1][1][DATA][26] ), .ZN(n1308) );
  AOI22_X1 U1515 ( .A1(n55), .A2(\cache[2][1][DATA][26] ), .B1(n237), .B2(
        \cache[3][1][DATA][26] ), .ZN(n1307) );
  AOI22_X1 U1516 ( .A1(n243), .A2(\cache[4][1][DATA][26] ), .B1(n241), .B2(
        \cache[5][1][DATA][26] ), .ZN(n1306) );
  AOI22_X1 U1517 ( .A1(n40), .A2(\cache[6][1][DATA][26] ), .B1(n245), .B2(
        \cache[7][1][DATA][26] ), .ZN(n1305) );
  AND4_X1 U1518 ( .A1(n1308), .A2(n1307), .A3(n1306), .A4(n1305), .ZN(n1327)
         );
  AOI22_X1 U1519 ( .A1(n233), .A2(\cache[0][0][DATA][26] ), .B1(n36), .B2(
        \cache[1][0][DATA][26] ), .ZN(n1312) );
  AOI22_X1 U1520 ( .A1(n240), .A2(\cache[2][0][DATA][26] ), .B1(n37), .B2(
        \cache[3][0][DATA][26] ), .ZN(n1311) );
  AOI22_X1 U1521 ( .A1(n56), .A2(\cache[4][0][DATA][26] ), .B1(n38), .B2(
        \cache[5][0][DATA][26] ), .ZN(n1310) );
  AOI22_X1 U1522 ( .A1(n40), .A2(\cache[6][0][DATA][26] ), .B1(n39), .B2(
        \cache[7][0][DATA][26] ), .ZN(n1309) );
  NAND4_X1 U1523 ( .A1(n1312), .A2(n1311), .A3(n1310), .A4(n1309), .ZN(n1319)
         );
  AOI22_X1 U1524 ( .A1(n233), .A2(\cache[0][2][DATA][26] ), .B1(n36), .B2(
        \cache[1][2][DATA][26] ), .ZN(n1316) );
  AOI22_X1 U1525 ( .A1(n55), .A2(\cache[2][2][DATA][26] ), .B1(n37), .B2(
        \cache[3][2][DATA][26] ), .ZN(n1315) );
  AOI22_X1 U1526 ( .A1(n56), .A2(\cache[4][2][DATA][26] ), .B1(n38), .B2(
        \cache[5][2][DATA][26] ), .ZN(n1314) );
  AOI22_X1 U1527 ( .A1(n40), .A2(\cache[6][2][DATA][26] ), .B1(n39), .B2(
        \cache[7][2][DATA][26] ), .ZN(n1313) );
  AND4_X1 U1528 ( .A1(n1316), .A2(n1315), .A3(n1314), .A4(n1313), .ZN(n1317)
         );
  AOI22_X1 U1529 ( .A1(n233), .A2(\cache[0][3][DATA][26] ), .B1(n36), .B2(
        \cache[1][3][DATA][26] ), .ZN(n1323) );
  AOI22_X1 U1530 ( .A1(n55), .A2(\cache[2][3][DATA][26] ), .B1(n37), .B2(
        \cache[3][3][DATA][26] ), .ZN(n1322) );
  AOI22_X1 U1531 ( .A1(n243), .A2(\cache[4][3][DATA][26] ), .B1(n38), .B2(
        \cache[5][3][DATA][26] ), .ZN(n1321) );
  AOI22_X1 U1532 ( .A1(n40), .A2(\cache[6][3][DATA][26] ), .B1(n39), .B2(
        \cache[7][3][DATA][26] ), .ZN(n1320) );
  NAND4_X1 U1533 ( .A1(n1323), .A2(n1322), .A3(n1321), .A4(n1320), .ZN(n1324)
         );
  AOI22_X1 U1534 ( .A1(n249), .A2(n1324), .B1(pc_in[28]), .B2(n91), .ZN(n1325)
         );
  OAI211_X1 U1535 ( .C1(n1327), .C2(n1584), .A(n1326), .B(n1325), .ZN(
        pc_out[28]) );
  AOI22_X1 U1536 ( .A1(n233), .A2(\cache[0][1][DATA][27] ), .B1(n231), .B2(
        \cache[1][1][DATA][27] ), .ZN(n1331) );
  AOI22_X1 U1537 ( .A1(n239), .A2(\cache[2][1][DATA][27] ), .B1(n237), .B2(
        \cache[3][1][DATA][27] ), .ZN(n1330) );
  AOI22_X1 U1538 ( .A1(n243), .A2(\cache[4][1][DATA][27] ), .B1(n241), .B2(
        \cache[5][1][DATA][27] ), .ZN(n1329) );
  AOI22_X1 U1539 ( .A1(n40), .A2(\cache[6][1][DATA][27] ), .B1(n245), .B2(
        \cache[7][1][DATA][27] ), .ZN(n1328) );
  AND4_X1 U1540 ( .A1(n1331), .A2(n1330), .A3(n1329), .A4(n1328), .ZN(n1350)
         );
  AOI22_X1 U1541 ( .A1(n235), .A2(\cache[0][0][DATA][27] ), .B1(n231), .B2(
        \cache[1][0][DATA][27] ), .ZN(n1335) );
  AOI22_X1 U1542 ( .A1(n239), .A2(\cache[2][0][DATA][27] ), .B1(n237), .B2(
        \cache[3][0][DATA][27] ), .ZN(n1334) );
  AOI22_X1 U1543 ( .A1(n243), .A2(\cache[4][0][DATA][27] ), .B1(n241), .B2(
        \cache[5][0][DATA][27] ), .ZN(n1333) );
  AOI22_X1 U1544 ( .A1(n40), .A2(\cache[6][0][DATA][27] ), .B1(n245), .B2(
        \cache[7][0][DATA][27] ), .ZN(n1332) );
  NAND4_X1 U1545 ( .A1(n1335), .A2(n1334), .A3(n1333), .A4(n1332), .ZN(n1342)
         );
  AOI22_X1 U1546 ( .A1(n235), .A2(\cache[0][2][DATA][27] ), .B1(n231), .B2(
        \cache[1][2][DATA][27] ), .ZN(n1339) );
  AOI22_X1 U1547 ( .A1(n239), .A2(\cache[2][2][DATA][27] ), .B1(n237), .B2(
        \cache[3][2][DATA][27] ), .ZN(n1338) );
  AOI22_X1 U1548 ( .A1(n243), .A2(\cache[4][2][DATA][27] ), .B1(n241), .B2(
        \cache[5][2][DATA][27] ), .ZN(n1337) );
  AOI22_X1 U1549 ( .A1(n40), .A2(\cache[6][2][DATA][27] ), .B1(n245), .B2(
        \cache[7][2][DATA][27] ), .ZN(n1336) );
  AND4_X1 U1550 ( .A1(n1339), .A2(n1338), .A3(n1337), .A4(n1336), .ZN(n1340)
         );
  AOI21_X1 U1551 ( .B1(n229), .B2(n1342), .A(n1341), .ZN(n1349) );
  AOI22_X1 U1552 ( .A1(n235), .A2(\cache[0][3][DATA][27] ), .B1(n231), .B2(
        \cache[1][3][DATA][27] ), .ZN(n1346) );
  AOI22_X1 U1553 ( .A1(n239), .A2(\cache[2][3][DATA][27] ), .B1(n237), .B2(
        \cache[3][3][DATA][27] ), .ZN(n1345) );
  AOI22_X1 U1554 ( .A1(n243), .A2(\cache[4][3][DATA][27] ), .B1(n241), .B2(
        \cache[5][3][DATA][27] ), .ZN(n1344) );
  AOI22_X1 U1555 ( .A1(n40), .A2(\cache[6][3][DATA][27] ), .B1(n245), .B2(
        \cache[7][3][DATA][27] ), .ZN(n1343) );
  NAND4_X1 U1556 ( .A1(n1346), .A2(n1345), .A3(n1344), .A4(n1343), .ZN(n1347)
         );
  AOI22_X1 U1557 ( .A1(n96), .A2(n1347), .B1(pc_in[29]), .B2(n91), .ZN(n1348)
         );
  AOI22_X1 U1558 ( .A1(n235), .A2(\cache[0][0][DATA][0] ), .B1(n231), .B2(
        \cache[1][0][DATA][0] ), .ZN(n1354) );
  AOI22_X1 U1559 ( .A1(n239), .A2(\cache[2][0][DATA][0] ), .B1(n237), .B2(
        \cache[3][0][DATA][0] ), .ZN(n1353) );
  AOI22_X1 U1560 ( .A1(n243), .A2(\cache[4][0][DATA][0] ), .B1(n241), .B2(
        \cache[5][0][DATA][0] ), .ZN(n1352) );
  AOI22_X1 U1561 ( .A1(n40), .A2(\cache[6][0][DATA][0] ), .B1(n245), .B2(
        \cache[7][0][DATA][0] ), .ZN(n1351) );
  NAND4_X1 U1562 ( .A1(n1354), .A2(n1353), .A3(n1352), .A4(n1351), .ZN(n1360)
         );
  AOI22_X1 U1563 ( .A1(n235), .A2(\cache[0][2][DATA][0] ), .B1(n231), .B2(
        \cache[1][2][DATA][0] ), .ZN(n1358) );
  AOI22_X1 U1564 ( .A1(n239), .A2(\cache[2][2][DATA][0] ), .B1(n237), .B2(
        \cache[3][2][DATA][0] ), .ZN(n1357) );
  AOI22_X1 U1565 ( .A1(n243), .A2(\cache[4][2][DATA][0] ), .B1(n241), .B2(
        \cache[5][2][DATA][0] ), .ZN(n1356) );
  AOI22_X1 U1566 ( .A1(n40), .A2(\cache[6][2][DATA][0] ), .B1(n245), .B2(
        \cache[7][2][DATA][0] ), .ZN(n1355) );
  AND4_X1 U1567 ( .A1(n1358), .A2(n1357), .A3(n1356), .A4(n1355), .ZN(n1359)
         );
  AOI22_X1 U1568 ( .A1(n235), .A2(\cache[0][1][DATA][0] ), .B1(n231), .B2(
        \cache[1][1][DATA][0] ), .ZN(n1364) );
  AOI22_X1 U1569 ( .A1(n239), .A2(\cache[2][1][DATA][0] ), .B1(n237), .B2(
        \cache[3][1][DATA][0] ), .ZN(n1363) );
  AOI22_X1 U1570 ( .A1(n243), .A2(\cache[4][1][DATA][0] ), .B1(n241), .B2(
        \cache[5][1][DATA][0] ), .ZN(n1362) );
  AOI22_X1 U1571 ( .A1(n40), .A2(\cache[6][1][DATA][0] ), .B1(n245), .B2(
        \cache[7][1][DATA][0] ), .ZN(n1361) );
  NAND4_X1 U1572 ( .A1(n1364), .A2(n1363), .A3(n1362), .A4(n1361), .ZN(n1370)
         );
  AOI22_X1 U1573 ( .A1(n235), .A2(\cache[0][3][DATA][0] ), .B1(n231), .B2(
        \cache[1][3][DATA][0] ), .ZN(n1368) );
  AOI22_X1 U1574 ( .A1(n239), .A2(\cache[2][3][DATA][0] ), .B1(n237), .B2(
        \cache[3][3][DATA][0] ), .ZN(n1367) );
  AOI22_X1 U1575 ( .A1(n243), .A2(\cache[4][3][DATA][0] ), .B1(n241), .B2(
        \cache[5][3][DATA][0] ), .ZN(n1366) );
  AOI22_X1 U1576 ( .A1(n40), .A2(\cache[6][3][DATA][0] ), .B1(n245), .B2(
        \cache[7][3][DATA][0] ), .ZN(n1365) );
  NAND4_X1 U1577 ( .A1(n1368), .A2(n1367), .A3(n1366), .A4(n1365), .ZN(n1369)
         );
  AOI22_X1 U1578 ( .A1(n235), .A2(\cache[0][1][DATA][28] ), .B1(n231), .B2(
        \cache[1][1][DATA][28] ), .ZN(n1376) );
  AOI22_X1 U1579 ( .A1(n239), .A2(\cache[2][1][DATA][28] ), .B1(n237), .B2(
        \cache[3][1][DATA][28] ), .ZN(n1375) );
  AOI22_X1 U1580 ( .A1(n243), .A2(\cache[4][1][DATA][28] ), .B1(n241), .B2(
        \cache[5][1][DATA][28] ), .ZN(n1374) );
  AOI22_X1 U1581 ( .A1(n40), .A2(\cache[6][1][DATA][28] ), .B1(n245), .B2(
        \cache[7][1][DATA][28] ), .ZN(n1373) );
  AND4_X1 U1582 ( .A1(n1376), .A2(n1375), .A3(n1374), .A4(n1373), .ZN(n1395)
         );
  AOI22_X1 U1583 ( .A1(n235), .A2(\cache[0][0][DATA][28] ), .B1(n231), .B2(
        \cache[1][0][DATA][28] ), .ZN(n1380) );
  AOI22_X1 U1584 ( .A1(n239), .A2(\cache[2][0][DATA][28] ), .B1(n237), .B2(
        \cache[3][0][DATA][28] ), .ZN(n1379) );
  AOI22_X1 U1585 ( .A1(n243), .A2(\cache[4][0][DATA][28] ), .B1(n241), .B2(
        \cache[5][0][DATA][28] ), .ZN(n1378) );
  AOI22_X1 U1586 ( .A1(n40), .A2(\cache[6][0][DATA][28] ), .B1(n245), .B2(
        \cache[7][0][DATA][28] ), .ZN(n1377) );
  NAND4_X1 U1587 ( .A1(n1380), .A2(n1379), .A3(n1378), .A4(n1377), .ZN(n1387)
         );
  AOI22_X1 U1588 ( .A1(n235), .A2(\cache[0][2][DATA][28] ), .B1(n231), .B2(
        \cache[1][2][DATA][28] ), .ZN(n1384) );
  AOI22_X1 U1589 ( .A1(n239), .A2(\cache[2][2][DATA][28] ), .B1(n237), .B2(
        \cache[3][2][DATA][28] ), .ZN(n1383) );
  AOI22_X1 U1590 ( .A1(n243), .A2(\cache[4][2][DATA][28] ), .B1(n241), .B2(
        \cache[5][2][DATA][28] ), .ZN(n1382) );
  AOI22_X1 U1591 ( .A1(n40), .A2(\cache[6][2][DATA][28] ), .B1(n245), .B2(
        \cache[7][2][DATA][28] ), .ZN(n1381) );
  AND4_X1 U1592 ( .A1(n1384), .A2(n1383), .A3(n1382), .A4(n1381), .ZN(n1385)
         );
  AOI22_X1 U1593 ( .A1(n235), .A2(\cache[0][3][DATA][28] ), .B1(n231), .B2(
        \cache[1][3][DATA][28] ), .ZN(n1391) );
  AOI22_X1 U1594 ( .A1(n55), .A2(\cache[2][3][DATA][28] ), .B1(n237), .B2(
        \cache[3][3][DATA][28] ), .ZN(n1390) );
  AOI22_X1 U1595 ( .A1(n56), .A2(\cache[4][3][DATA][28] ), .B1(n241), .B2(
        \cache[5][3][DATA][28] ), .ZN(n1389) );
  AOI22_X1 U1596 ( .A1(n40), .A2(\cache[6][3][DATA][28] ), .B1(n245), .B2(
        \cache[7][3][DATA][28] ), .ZN(n1388) );
  NAND4_X1 U1597 ( .A1(n1391), .A2(n1390), .A3(n1389), .A4(n1388), .ZN(n1392)
         );
  AOI22_X1 U1598 ( .A1(n249), .A2(n1392), .B1(pc_in[30]), .B2(n91), .ZN(n1393)
         );
  OAI211_X1 U1599 ( .C1(n1395), .C2(n1584), .A(n1394), .B(n1393), .ZN(
        pc_out[30]) );
  AOI22_X1 U1600 ( .A1(n233), .A2(\cache[0][1][DATA][29] ), .B1(n231), .B2(
        \cache[1][1][DATA][29] ), .ZN(n1399) );
  AOI22_X1 U1601 ( .A1(n55), .A2(\cache[2][1][DATA][29] ), .B1(n237), .B2(
        \cache[3][1][DATA][29] ), .ZN(n1398) );
  AOI22_X1 U1602 ( .A1(n56), .A2(\cache[4][1][DATA][29] ), .B1(n241), .B2(
        \cache[5][1][DATA][29] ), .ZN(n1397) );
  AOI22_X1 U1603 ( .A1(n40), .A2(\cache[6][1][DATA][29] ), .B1(n245), .B2(
        \cache[7][1][DATA][29] ), .ZN(n1396) );
  AND4_X1 U1604 ( .A1(n1399), .A2(n1398), .A3(n1397), .A4(n1396), .ZN(n1416)
         );
  AOI22_X1 U1605 ( .A1(n233), .A2(\cache[0][0][DATA][29] ), .B1(n231), .B2(
        \cache[1][0][DATA][29] ), .ZN(n1403) );
  AOI22_X1 U1606 ( .A1(n55), .A2(\cache[2][0][DATA][29] ), .B1(n237), .B2(
        \cache[3][0][DATA][29] ), .ZN(n1402) );
  AOI22_X1 U1607 ( .A1(n56), .A2(\cache[4][0][DATA][29] ), .B1(n241), .B2(
        \cache[5][0][DATA][29] ), .ZN(n1401) );
  AOI22_X1 U1608 ( .A1(n40), .A2(\cache[6][0][DATA][29] ), .B1(n245), .B2(
        \cache[7][0][DATA][29] ), .ZN(n1400) );
  NAND4_X1 U1609 ( .A1(n1403), .A2(n1402), .A3(n1401), .A4(n1400), .ZN(n1410)
         );
  AOI22_X1 U1610 ( .A1(n233), .A2(\cache[0][2][DATA][29] ), .B1(n231), .B2(
        \cache[1][2][DATA][29] ), .ZN(n1407) );
  AOI22_X1 U1611 ( .A1(n55), .A2(\cache[2][2][DATA][29] ), .B1(n237), .B2(
        \cache[3][2][DATA][29] ), .ZN(n1406) );
  AOI22_X1 U1612 ( .A1(n56), .A2(\cache[4][2][DATA][29] ), .B1(n241), .B2(
        \cache[5][2][DATA][29] ), .ZN(n1405) );
  AOI22_X1 U1613 ( .A1(n40), .A2(\cache[6][2][DATA][29] ), .B1(n245), .B2(
        \cache[7][2][DATA][29] ), .ZN(n1404) );
  AND4_X1 U1614 ( .A1(n1407), .A2(n1406), .A3(n1405), .A4(n1404), .ZN(n1408)
         );
  AOI22_X1 U1615 ( .A1(n233), .A2(\cache[0][3][DATA][29] ), .B1(n231), .B2(
        \cache[1][3][DATA][29] ), .ZN(n1414) );
  AOI22_X1 U1616 ( .A1(n55), .A2(\cache[2][3][DATA][29] ), .B1(n237), .B2(
        \cache[3][3][DATA][29] ), .ZN(n1413) );
  AOI22_X1 U1617 ( .A1(n56), .A2(\cache[4][3][DATA][29] ), .B1(n241), .B2(
        \cache[5][3][DATA][29] ), .ZN(n1412) );
  AOI22_X1 U1618 ( .A1(n40), .A2(\cache[6][3][DATA][29] ), .B1(n245), .B2(
        \cache[7][3][DATA][29] ), .ZN(n1411) );
  NAND4_X1 U1619 ( .A1(n1414), .A2(n1413), .A3(n1412), .A4(n1411), .ZN(n1415)
         );
  AOI22_X1 U1620 ( .A1(n233), .A2(\cache[0][1][DATA][1] ), .B1(n231), .B2(
        \cache[1][1][DATA][1] ), .ZN(n1420) );
  AOI22_X1 U1621 ( .A1(n55), .A2(\cache[2][1][DATA][1] ), .B1(n237), .B2(
        \cache[3][1][DATA][1] ), .ZN(n1419) );
  AOI22_X1 U1622 ( .A1(n56), .A2(\cache[4][1][DATA][1] ), .B1(n241), .B2(
        \cache[5][1][DATA][1] ), .ZN(n1418) );
  AOI22_X1 U1623 ( .A1(n40), .A2(\cache[6][1][DATA][1] ), .B1(n245), .B2(
        \cache[7][1][DATA][1] ), .ZN(n1417) );
  AND4_X1 U1624 ( .A1(n1420), .A2(n1419), .A3(n1418), .A4(n1417), .ZN(n1439)
         );
  AOI22_X1 U1625 ( .A1(n233), .A2(\cache[0][0][DATA][1] ), .B1(n231), .B2(
        \cache[1][0][DATA][1] ), .ZN(n1424) );
  AOI22_X1 U1626 ( .A1(n55), .A2(\cache[2][0][DATA][1] ), .B1(n237), .B2(
        \cache[3][0][DATA][1] ), .ZN(n1423) );
  AOI22_X1 U1627 ( .A1(n56), .A2(\cache[4][0][DATA][1] ), .B1(n241), .B2(
        \cache[5][0][DATA][1] ), .ZN(n1422) );
  AOI22_X1 U1628 ( .A1(n40), .A2(\cache[6][0][DATA][1] ), .B1(n245), .B2(
        \cache[7][0][DATA][1] ), .ZN(n1421) );
  NAND4_X1 U1629 ( .A1(n1424), .A2(n1423), .A3(n1422), .A4(n1421), .ZN(n1431)
         );
  AOI22_X1 U1630 ( .A1(n233), .A2(\cache[0][2][DATA][1] ), .B1(n231), .B2(
        \cache[1][2][DATA][1] ), .ZN(n1428) );
  AOI22_X1 U1631 ( .A1(n55), .A2(\cache[2][2][DATA][1] ), .B1(n237), .B2(
        \cache[3][2][DATA][1] ), .ZN(n1427) );
  AOI22_X1 U1632 ( .A1(n56), .A2(\cache[4][2][DATA][1] ), .B1(n241), .B2(
        \cache[5][2][DATA][1] ), .ZN(n1426) );
  AOI22_X1 U1633 ( .A1(n40), .A2(\cache[6][2][DATA][1] ), .B1(n245), .B2(
        \cache[7][2][DATA][1] ), .ZN(n1425) );
  AND4_X1 U1634 ( .A1(n1428), .A2(n1427), .A3(n1426), .A4(n1425), .ZN(n1429)
         );
  AOI21_X1 U1635 ( .B1(n230), .B2(n1431), .A(n1430), .ZN(n1438) );
  AOI22_X1 U1636 ( .A1(n233), .A2(\cache[0][3][DATA][1] ), .B1(n231), .B2(
        \cache[1][3][DATA][1] ), .ZN(n1435) );
  AOI22_X1 U1637 ( .A1(n55), .A2(\cache[2][3][DATA][1] ), .B1(n237), .B2(
        \cache[3][3][DATA][1] ), .ZN(n1434) );
  AOI22_X1 U1638 ( .A1(n56), .A2(\cache[4][3][DATA][1] ), .B1(n241), .B2(
        \cache[5][3][DATA][1] ), .ZN(n1433) );
  AOI22_X1 U1639 ( .A1(n40), .A2(\cache[6][3][DATA][1] ), .B1(n245), .B2(
        \cache[7][3][DATA][1] ), .ZN(n1432) );
  NAND4_X1 U1640 ( .A1(n1435), .A2(n1434), .A3(n1433), .A4(n1432), .ZN(n1436)
         );
  AOI22_X1 U1641 ( .A1(n249), .A2(n1436), .B1(pc_in[3]), .B2(n91), .ZN(n1437)
         );
  AOI22_X1 U1642 ( .A1(n233), .A2(\cache[0][1][DATA][2] ), .B1(n231), .B2(
        \cache[1][1][DATA][2] ), .ZN(n1443) );
  AOI22_X1 U1643 ( .A1(n55), .A2(\cache[2][1][DATA][2] ), .B1(n237), .B2(
        \cache[3][1][DATA][2] ), .ZN(n1442) );
  AOI22_X1 U1644 ( .A1(n56), .A2(\cache[4][1][DATA][2] ), .B1(n241), .B2(
        \cache[5][1][DATA][2] ), .ZN(n1441) );
  AOI22_X1 U1645 ( .A1(n40), .A2(\cache[6][1][DATA][2] ), .B1(n245), .B2(
        \cache[7][1][DATA][2] ), .ZN(n1440) );
  AND4_X1 U1646 ( .A1(n1443), .A2(n1442), .A3(n1441), .A4(n1440), .ZN(n1460)
         );
  AOI22_X1 U1647 ( .A1(n233), .A2(\cache[0][0][DATA][2] ), .B1(n231), .B2(
        \cache[1][0][DATA][2] ), .ZN(n1447) );
  AOI22_X1 U1648 ( .A1(n55), .A2(\cache[2][0][DATA][2] ), .B1(n237), .B2(
        \cache[3][0][DATA][2] ), .ZN(n1446) );
  AOI22_X1 U1649 ( .A1(n56), .A2(\cache[4][0][DATA][2] ), .B1(n241), .B2(
        \cache[5][0][DATA][2] ), .ZN(n1445) );
  AOI22_X1 U1650 ( .A1(n40), .A2(\cache[6][0][DATA][2] ), .B1(n245), .B2(
        \cache[7][0][DATA][2] ), .ZN(n1444) );
  NAND4_X1 U1651 ( .A1(n1447), .A2(n1446), .A3(n1445), .A4(n1444), .ZN(n1454)
         );
  AOI22_X1 U1652 ( .A1(n233), .A2(\cache[0][2][DATA][2] ), .B1(n231), .B2(
        \cache[1][2][DATA][2] ), .ZN(n1451) );
  AOI22_X1 U1653 ( .A1(n239), .A2(\cache[2][2][DATA][2] ), .B1(n237), .B2(
        \cache[3][2][DATA][2] ), .ZN(n1450) );
  AOI22_X1 U1654 ( .A1(n243), .A2(\cache[4][2][DATA][2] ), .B1(n241), .B2(
        \cache[5][2][DATA][2] ), .ZN(n1449) );
  AOI22_X1 U1655 ( .A1(n40), .A2(\cache[6][2][DATA][2] ), .B1(n245), .B2(
        \cache[7][2][DATA][2] ), .ZN(n1448) );
  AND4_X1 U1656 ( .A1(n1451), .A2(n1450), .A3(n1449), .A4(n1448), .ZN(n1452)
         );
  AOI22_X1 U1657 ( .A1(n57), .A2(\cache[0][3][DATA][2] ), .B1(n231), .B2(
        \cache[1][3][DATA][2] ), .ZN(n1458) );
  AOI22_X1 U1658 ( .A1(n239), .A2(\cache[2][3][DATA][2] ), .B1(n237), .B2(
        \cache[3][3][DATA][2] ), .ZN(n1457) );
  AOI22_X1 U1659 ( .A1(n243), .A2(\cache[4][3][DATA][2] ), .B1(n241), .B2(
        \cache[5][3][DATA][2] ), .ZN(n1456) );
  AOI22_X1 U1660 ( .A1(n40), .A2(\cache[6][3][DATA][2] ), .B1(n245), .B2(
        \cache[7][3][DATA][2] ), .ZN(n1455) );
  NAND4_X1 U1661 ( .A1(n1458), .A2(n1457), .A3(n1456), .A4(n1455), .ZN(n1459)
         );
  AOI22_X1 U1662 ( .A1(n57), .A2(\cache[0][1][DATA][3] ), .B1(n231), .B2(
        \cache[1][1][DATA][3] ), .ZN(n1464) );
  AOI22_X1 U1663 ( .A1(n239), .A2(\cache[2][1][DATA][3] ), .B1(n237), .B2(
        \cache[3][1][DATA][3] ), .ZN(n1463) );
  AOI22_X1 U1664 ( .A1(n243), .A2(\cache[4][1][DATA][3] ), .B1(n241), .B2(
        \cache[5][1][DATA][3] ), .ZN(n1462) );
  AOI22_X1 U1665 ( .A1(n40), .A2(\cache[6][1][DATA][3] ), .B1(n245), .B2(
        \cache[7][1][DATA][3] ), .ZN(n1461) );
  AND4_X1 U1666 ( .A1(n1464), .A2(n1463), .A3(n1462), .A4(n1461), .ZN(n1481)
         );
  AOI22_X1 U1667 ( .A1(n57), .A2(\cache[0][0][DATA][3] ), .B1(n231), .B2(
        \cache[1][0][DATA][3] ), .ZN(n1468) );
  AOI22_X1 U1668 ( .A1(n239), .A2(\cache[2][0][DATA][3] ), .B1(n237), .B2(
        \cache[3][0][DATA][3] ), .ZN(n1467) );
  AOI22_X1 U1669 ( .A1(n243), .A2(\cache[4][0][DATA][3] ), .B1(n241), .B2(
        \cache[5][0][DATA][3] ), .ZN(n1466) );
  AOI22_X1 U1670 ( .A1(n40), .A2(\cache[6][0][DATA][3] ), .B1(n245), .B2(
        \cache[7][0][DATA][3] ), .ZN(n1465) );
  NAND4_X1 U1671 ( .A1(n1468), .A2(n1467), .A3(n1466), .A4(n1465), .ZN(n1475)
         );
  AOI22_X1 U1672 ( .A1(n57), .A2(\cache[0][2][DATA][3] ), .B1(n231), .B2(
        \cache[1][2][DATA][3] ), .ZN(n1472) );
  AOI22_X1 U1673 ( .A1(n239), .A2(\cache[2][2][DATA][3] ), .B1(n237), .B2(
        \cache[3][2][DATA][3] ), .ZN(n1471) );
  AOI22_X1 U1674 ( .A1(n243), .A2(\cache[4][2][DATA][3] ), .B1(n241), .B2(
        \cache[5][2][DATA][3] ), .ZN(n1470) );
  AOI22_X1 U1675 ( .A1(n40), .A2(\cache[6][2][DATA][3] ), .B1(n245), .B2(
        \cache[7][2][DATA][3] ), .ZN(n1469) );
  AND4_X1 U1676 ( .A1(n1472), .A2(n1471), .A3(n1470), .A4(n1469), .ZN(n1473)
         );
  AOI22_X1 U1677 ( .A1(n57), .A2(\cache[0][3][DATA][3] ), .B1(n231), .B2(
        \cache[1][3][DATA][3] ), .ZN(n1479) );
  AOI22_X1 U1678 ( .A1(n239), .A2(\cache[2][3][DATA][3] ), .B1(n237), .B2(
        \cache[3][3][DATA][3] ), .ZN(n1478) );
  AOI22_X1 U1679 ( .A1(n243), .A2(\cache[4][3][DATA][3] ), .B1(n241), .B2(
        \cache[5][3][DATA][3] ), .ZN(n1477) );
  AOI22_X1 U1680 ( .A1(n40), .A2(\cache[6][3][DATA][3] ), .B1(n245), .B2(
        \cache[7][3][DATA][3] ), .ZN(n1476) );
  NAND4_X1 U1681 ( .A1(n1479), .A2(n1478), .A3(n1477), .A4(n1476), .ZN(n1480)
         );
  AOI22_X1 U1682 ( .A1(n57), .A2(\cache[0][1][DATA][4] ), .B1(n231), .B2(
        \cache[1][1][DATA][4] ), .ZN(n1485) );
  AOI22_X1 U1683 ( .A1(n239), .A2(\cache[2][1][DATA][4] ), .B1(n237), .B2(
        \cache[3][1][DATA][4] ), .ZN(n1484) );
  AOI22_X1 U1684 ( .A1(n243), .A2(\cache[4][1][DATA][4] ), .B1(n241), .B2(
        \cache[5][1][DATA][4] ), .ZN(n1483) );
  AOI22_X1 U1685 ( .A1(n40), .A2(\cache[6][1][DATA][4] ), .B1(n245), .B2(
        \cache[7][1][DATA][4] ), .ZN(n1482) );
  AND4_X1 U1686 ( .A1(n1485), .A2(n1484), .A3(n1483), .A4(n1482), .ZN(n1504)
         );
  AOI22_X1 U1687 ( .A1(n57), .A2(\cache[0][0][DATA][4] ), .B1(n231), .B2(
        \cache[1][0][DATA][4] ), .ZN(n1489) );
  AOI22_X1 U1688 ( .A1(n239), .A2(\cache[2][0][DATA][4] ), .B1(n237), .B2(
        \cache[3][0][DATA][4] ), .ZN(n1488) );
  AOI22_X1 U1689 ( .A1(n243), .A2(\cache[4][0][DATA][4] ), .B1(n241), .B2(
        \cache[5][0][DATA][4] ), .ZN(n1487) );
  AOI22_X1 U1690 ( .A1(n40), .A2(\cache[6][0][DATA][4] ), .B1(n245), .B2(
        \cache[7][0][DATA][4] ), .ZN(n1486) );
  NAND4_X1 U1691 ( .A1(n1489), .A2(n1488), .A3(n1487), .A4(n1486), .ZN(n1496)
         );
  AOI22_X1 U1692 ( .A1(n233), .A2(\cache[0][2][DATA][4] ), .B1(n36), .B2(
        \cache[1][2][DATA][4] ), .ZN(n1493) );
  AOI22_X1 U1693 ( .A1(n239), .A2(\cache[2][2][DATA][4] ), .B1(n37), .B2(
        \cache[3][2][DATA][4] ), .ZN(n1492) );
  AOI22_X1 U1694 ( .A1(n243), .A2(\cache[4][2][DATA][4] ), .B1(n38), .B2(
        \cache[5][2][DATA][4] ), .ZN(n1491) );
  AOI22_X1 U1695 ( .A1(n40), .A2(\cache[6][2][DATA][4] ), .B1(n39), .B2(
        \cache[7][2][DATA][4] ), .ZN(n1490) );
  AND4_X1 U1696 ( .A1(n1493), .A2(n1492), .A3(n1491), .A4(n1490), .ZN(n1494)
         );
  AOI21_X1 U1697 ( .B1(n230), .B2(n1496), .A(n1495), .ZN(n1503) );
  AOI22_X1 U1698 ( .A1(n57), .A2(\cache[0][3][DATA][4] ), .B1(n231), .B2(
        \cache[1][3][DATA][4] ), .ZN(n1500) );
  AOI22_X1 U1699 ( .A1(n239), .A2(\cache[2][3][DATA][4] ), .B1(n237), .B2(
        \cache[3][3][DATA][4] ), .ZN(n1499) );
  AOI22_X1 U1700 ( .A1(n243), .A2(\cache[4][3][DATA][4] ), .B1(n241), .B2(
        \cache[5][3][DATA][4] ), .ZN(n1498) );
  AOI22_X1 U1701 ( .A1(n40), .A2(\cache[6][3][DATA][4] ), .B1(n245), .B2(
        \cache[7][3][DATA][4] ), .ZN(n1497) );
  NAND4_X1 U1702 ( .A1(n1500), .A2(n1499), .A3(n1498), .A4(n1497), .ZN(n1501)
         );
  AOI22_X1 U1703 ( .A1(n96), .A2(n1501), .B1(pc_in[6]), .B2(n93), .ZN(n1502)
         );
  AOI22_X1 U1704 ( .A1(n233), .A2(\cache[0][1][DATA][5] ), .B1(n36), .B2(
        \cache[1][1][DATA][5] ), .ZN(n1508) );
  AOI22_X1 U1705 ( .A1(n239), .A2(\cache[2][1][DATA][5] ), .B1(n37), .B2(
        \cache[3][1][DATA][5] ), .ZN(n1507) );
  AOI22_X1 U1706 ( .A1(n243), .A2(\cache[4][1][DATA][5] ), .B1(n38), .B2(
        \cache[5][1][DATA][5] ), .ZN(n1506) );
  AOI22_X1 U1707 ( .A1(n40), .A2(\cache[6][1][DATA][5] ), .B1(n39), .B2(
        \cache[7][1][DATA][5] ), .ZN(n1505) );
  AND4_X1 U1708 ( .A1(n1508), .A2(n1507), .A3(n1506), .A4(n1505), .ZN(n1527)
         );
  AOI22_X1 U1709 ( .A1(n233), .A2(\cache[0][0][DATA][5] ), .B1(n36), .B2(
        \cache[1][0][DATA][5] ), .ZN(n1512) );
  AOI22_X1 U1710 ( .A1(n240), .A2(\cache[2][0][DATA][5] ), .B1(n37), .B2(
        \cache[3][0][DATA][5] ), .ZN(n1511) );
  AOI22_X1 U1711 ( .A1(n244), .A2(\cache[4][0][DATA][5] ), .B1(n38), .B2(
        \cache[5][0][DATA][5] ), .ZN(n1510) );
  AOI22_X1 U1712 ( .A1(n40), .A2(\cache[6][0][DATA][5] ), .B1(n39), .B2(
        \cache[7][0][DATA][5] ), .ZN(n1509) );
  NAND4_X1 U1713 ( .A1(n1512), .A2(n1511), .A3(n1510), .A4(n1509), .ZN(n1519)
         );
  AOI22_X1 U1714 ( .A1(n57), .A2(\cache[0][2][DATA][5] ), .B1(n231), .B2(
        \cache[1][2][DATA][5] ), .ZN(n1516) );
  AOI22_X1 U1715 ( .A1(n240), .A2(\cache[2][2][DATA][5] ), .B1(n237), .B2(
        \cache[3][2][DATA][5] ), .ZN(n1515) );
  AOI22_X1 U1716 ( .A1(n244), .A2(\cache[4][2][DATA][5] ), .B1(n241), .B2(
        \cache[5][2][DATA][5] ), .ZN(n1514) );
  AOI22_X1 U1717 ( .A1(n40), .A2(\cache[6][2][DATA][5] ), .B1(n245), .B2(
        \cache[7][2][DATA][5] ), .ZN(n1513) );
  AND4_X1 U1718 ( .A1(n1516), .A2(n1515), .A3(n1514), .A4(n1513), .ZN(n1517)
         );
  AOI21_X1 U1719 ( .B1(n25), .B2(n1519), .A(n1518), .ZN(n1526) );
  AOI22_X1 U1720 ( .A1(n235), .A2(\cache[0][3][DATA][5] ), .B1(n36), .B2(
        \cache[1][3][DATA][5] ), .ZN(n1523) );
  AOI22_X1 U1721 ( .A1(n240), .A2(\cache[2][3][DATA][5] ), .B1(n37), .B2(
        \cache[3][3][DATA][5] ), .ZN(n1522) );
  AOI22_X1 U1722 ( .A1(n244), .A2(\cache[4][3][DATA][5] ), .B1(n38), .B2(
        \cache[5][3][DATA][5] ), .ZN(n1521) );
  AOI22_X1 U1723 ( .A1(n40), .A2(\cache[6][3][DATA][5] ), .B1(n39), .B2(
        \cache[7][3][DATA][5] ), .ZN(n1520) );
  NAND4_X1 U1724 ( .A1(n1523), .A2(n1522), .A3(n1521), .A4(n1520), .ZN(n1524)
         );
  AOI22_X1 U1725 ( .A1(n249), .A2(n1524), .B1(pc_in[7]), .B2(n93), .ZN(n1525)
         );
  AOI22_X1 U1726 ( .A1(n235), .A2(\cache[0][1][DATA][6] ), .B1(n36), .B2(
        \cache[1][1][DATA][6] ), .ZN(n1531) );
  AOI22_X1 U1727 ( .A1(n239), .A2(\cache[2][1][DATA][6] ), .B1(n37), .B2(
        \cache[3][1][DATA][6] ), .ZN(n1530) );
  AOI22_X1 U1728 ( .A1(n243), .A2(\cache[4][1][DATA][6] ), .B1(n38), .B2(
        \cache[5][1][DATA][6] ), .ZN(n1529) );
  AOI22_X1 U1729 ( .A1(n40), .A2(\cache[6][1][DATA][6] ), .B1(n39), .B2(
        \cache[7][1][DATA][6] ), .ZN(n1528) );
  AND4_X1 U1730 ( .A1(n1531), .A2(n1530), .A3(n1529), .A4(n1528), .ZN(n1550)
         );
  AOI22_X1 U1731 ( .A1(n57), .A2(\cache[0][0][DATA][6] ), .B1(n231), .B2(
        \cache[1][0][DATA][6] ), .ZN(n1535) );
  AOI22_X1 U1732 ( .A1(n240), .A2(\cache[2][0][DATA][6] ), .B1(n237), .B2(
        \cache[3][0][DATA][6] ), .ZN(n1534) );
  AOI22_X1 U1733 ( .A1(n244), .A2(\cache[4][0][DATA][6] ), .B1(n241), .B2(
        \cache[5][0][DATA][6] ), .ZN(n1533) );
  AOI22_X1 U1734 ( .A1(n40), .A2(\cache[6][0][DATA][6] ), .B1(n245), .B2(
        \cache[7][0][DATA][6] ), .ZN(n1532) );
  NAND4_X1 U1735 ( .A1(n1535), .A2(n1534), .A3(n1533), .A4(n1532), .ZN(n1542)
         );
  AOI22_X1 U1736 ( .A1(n235), .A2(\cache[0][2][DATA][6] ), .B1(n36), .B2(
        \cache[1][2][DATA][6] ), .ZN(n1539) );
  AOI22_X1 U1737 ( .A1(n240), .A2(\cache[2][2][DATA][6] ), .B1(n37), .B2(
        \cache[3][2][DATA][6] ), .ZN(n1538) );
  AOI22_X1 U1738 ( .A1(n244), .A2(\cache[4][2][DATA][6] ), .B1(n38), .B2(
        \cache[5][2][DATA][6] ), .ZN(n1537) );
  AOI22_X1 U1739 ( .A1(n40), .A2(\cache[6][2][DATA][6] ), .B1(n39), .B2(
        \cache[7][2][DATA][6] ), .ZN(n1536) );
  AND4_X1 U1740 ( .A1(n1539), .A2(n1538), .A3(n1537), .A4(n1536), .ZN(n1540)
         );
  AOI21_X1 U1741 ( .B1(n229), .B2(n1542), .A(n1541), .ZN(n1549) );
  AOI22_X1 U1742 ( .A1(n233), .A2(\cache[0][3][DATA][6] ), .B1(n36), .B2(
        \cache[1][3][DATA][6] ), .ZN(n1546) );
  AOI22_X1 U1743 ( .A1(n240), .A2(\cache[2][3][DATA][6] ), .B1(n37), .B2(
        \cache[3][3][DATA][6] ), .ZN(n1545) );
  AOI22_X1 U1744 ( .A1(n244), .A2(\cache[4][3][DATA][6] ), .B1(n38), .B2(
        \cache[5][3][DATA][6] ), .ZN(n1544) );
  AOI22_X1 U1745 ( .A1(n40), .A2(\cache[6][3][DATA][6] ), .B1(n39), .B2(
        \cache[7][3][DATA][6] ), .ZN(n1543) );
  NAND4_X1 U1746 ( .A1(n1546), .A2(n1545), .A3(n1544), .A4(n1543), .ZN(n1547)
         );
  AOI22_X1 U1747 ( .A1(n96), .A2(n1547), .B1(pc_in[8]), .B2(n93), .ZN(n1548)
         );
  AOI22_X1 U1748 ( .A1(n235), .A2(\cache[0][1][DATA][7] ), .B1(n36), .B2(
        \cache[1][1][DATA][7] ), .ZN(n1554) );
  AOI22_X1 U1749 ( .A1(n239), .A2(\cache[2][1][DATA][7] ), .B1(n37), .B2(
        \cache[3][1][DATA][7] ), .ZN(n1553) );
  AOI22_X1 U1750 ( .A1(n243), .A2(\cache[4][1][DATA][7] ), .B1(n38), .B2(
        \cache[5][1][DATA][7] ), .ZN(n1552) );
  AOI22_X1 U1751 ( .A1(n40), .A2(\cache[6][1][DATA][7] ), .B1(n39), .B2(
        \cache[7][1][DATA][7] ), .ZN(n1551) );
  AND4_X1 U1752 ( .A1(n1554), .A2(n1553), .A3(n1552), .A4(n1551), .ZN(n1585)
         );
  AOI22_X1 U1753 ( .A1(n57), .A2(\cache[0][0][DATA][7] ), .B1(n231), .B2(
        \cache[1][0][DATA][7] ), .ZN(n1558) );
  AOI22_X1 U1754 ( .A1(n240), .A2(\cache[2][0][DATA][7] ), .B1(n237), .B2(
        \cache[3][0][DATA][7] ), .ZN(n1557) );
  AOI22_X1 U1755 ( .A1(n244), .A2(\cache[4][0][DATA][7] ), .B1(n241), .B2(
        \cache[5][0][DATA][7] ), .ZN(n1556) );
  AOI22_X1 U1756 ( .A1(n40), .A2(\cache[6][0][DATA][7] ), .B1(n245), .B2(
        \cache[7][0][DATA][7] ), .ZN(n1555) );
  NAND4_X1 U1757 ( .A1(n1558), .A2(n1557), .A3(n1556), .A4(n1555), .ZN(n1566)
         );
  AOI22_X1 U1758 ( .A1(n233), .A2(\cache[0][2][DATA][7] ), .B1(n36), .B2(
        \cache[1][2][DATA][7] ), .ZN(n1562) );
  AOI22_X1 U1759 ( .A1(n240), .A2(\cache[2][2][DATA][7] ), .B1(n37), .B2(
        \cache[3][2][DATA][7] ), .ZN(n1561) );
  AOI22_X1 U1760 ( .A1(n244), .A2(\cache[4][2][DATA][7] ), .B1(n38), .B2(
        \cache[5][2][DATA][7] ), .ZN(n1560) );
  AOI22_X1 U1761 ( .A1(n40), .A2(\cache[6][2][DATA][7] ), .B1(n39), .B2(
        \cache[7][2][DATA][7] ), .ZN(n1559) );
  AND4_X1 U1762 ( .A1(n1562), .A2(n1561), .A3(n1560), .A4(n1559), .ZN(n1564)
         );
  AOI21_X1 U1763 ( .B1(n229), .B2(n1566), .A(n1565), .ZN(n1583) );
  AOI22_X1 U1764 ( .A1(n236), .A2(\cache[0][3][DATA][7] ), .B1(n36), .B2(
        \cache[1][3][DATA][7] ), .ZN(n1579) );
  AOI22_X1 U1765 ( .A1(n239), .A2(\cache[2][3][DATA][7] ), .B1(n37), .B2(
        \cache[3][3][DATA][7] ), .ZN(n1578) );
  AOI22_X1 U1766 ( .A1(n243), .A2(\cache[4][3][DATA][7] ), .B1(n38), .B2(
        \cache[5][3][DATA][7] ), .ZN(n1577) );
  AOI22_X1 U1767 ( .A1(n40), .A2(\cache[6][3][DATA][7] ), .B1(n246), .B2(
        \cache[7][3][DATA][7] ), .ZN(n1576) );
  NAND4_X1 U1768 ( .A1(n1579), .A2(n1578), .A3(n1577), .A4(n1576), .ZN(n1580)
         );
  AOI22_X1 U1769 ( .A1(n96), .A2(n1580), .B1(pc_in[9]), .B2(n93), .ZN(n1582)
         );
endmodule


module SNPS_CLOCK_GATE_HIGH_reg_N32_12 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18782, net18784, net18786, net18787, net18790, net18793;
  assign net18782 = EN;
  assign net18784 = CLK;
  assign ENCLK = net18786;
  assign net18793 = TE;

  DLL_X1 latch ( .D(net18787), .GN(net18784), .Q(net18790) );
  AND2_X1 main_gate ( .A1(net18790), .A2(net18784), .ZN(net18786) );
  OR2_X1 test_or ( .A1(net18782), .A2(net18793), .ZN(net18787) );
endmodule


module reg_N32_12 ( Q, EN, CLK, RST, \D[31] , \D[30] , \D[29] , \D[28] , 
        \D[27] , \D[26] , \D[25] , \D[24] , \D[23] , \D[22] , \D[21] , \D[20] , 
        \D[19] , \D[18] , \D[17] , \D[16] , \D[15] , \D[14] , \D[13] , \D[12] , 
        \D[11] , \D[10] , \D[9] , \D[8] , \D[7] , \D[6] , \D[5] , \D[4] , 
        \D[3] , \D[2]_BAR , \D[1] , \D[0]  );
  output [31:0] Q;
  input EN, CLK, RST, \D[31] , \D[30] , \D[29] , \D[28] , \D[27] , \D[26] ,
         \D[25] , \D[24] , \D[23] , \D[22] , \D[21] , \D[20] , \D[19] ,
         \D[18] , \D[17] , \D[16] , \D[15] , \D[14] , \D[13] , \D[12] ,
         \D[11] , \D[10] , \D[9] , \D[8] , \D[7] , \D[6] , \D[5] , \D[4] ,
         \D[3] , \D[2]_BAR , \D[1] , \D[0] ;
  wire   net18798, n1;
  wire   [31:0] D;
  assign D[2] = \D[2]_BAR ;

  SNPS_CLOCK_GATE_HIGH_reg_N32_12 clk_gate_Q_reg ( .CLK(CLK), .EN(EN), .ENCLK(
        net18798), .TE(1'b0) );
  DFFR_X1 \Q_reg[31]  ( .D(D[31]), .CK(net18798), .RN(RST), .Q(Q[31]) );
  DFFR_X1 \Q_reg[30]  ( .D(D[30]), .CK(net18798), .RN(RST), .Q(Q[30]) );
  DFFR_X1 \Q_reg[29]  ( .D(D[29]), .CK(net18798), .RN(RST), .Q(Q[29]) );
  DFFR_X1 \Q_reg[28]  ( .D(D[28]), .CK(net18798), .RN(RST), .Q(Q[28]) );
  DFFR_X1 \Q_reg[27]  ( .D(D[27]), .CK(net18798), .RN(RST), .Q(Q[27]) );
  DFFR_X1 \Q_reg[26]  ( .D(D[26]), .CK(net18798), .RN(RST), .Q(Q[26]) );
  DFFR_X1 \Q_reg[25]  ( .D(D[25]), .CK(net18798), .RN(RST), .Q(Q[25]) );
  DFFR_X1 \Q_reg[24]  ( .D(D[24]), .CK(net18798), .RN(RST), .Q(Q[24]) );
  DFFR_X1 \Q_reg[23]  ( .D(D[23]), .CK(net18798), .RN(RST), .Q(Q[23]) );
  DFFR_X1 \Q_reg[22]  ( .D(D[22]), .CK(net18798), .RN(RST), .Q(Q[22]) );
  DFFR_X1 \Q_reg[21]  ( .D(D[21]), .CK(net18798), .RN(RST), .Q(Q[21]) );
  DFFR_X1 \Q_reg[20]  ( .D(D[20]), .CK(net18798), .RN(RST), .Q(Q[20]) );
  DFFR_X1 \Q_reg[19]  ( .D(D[19]), .CK(net18798), .RN(RST), .Q(Q[19]) );
  DFFR_X1 \Q_reg[18]  ( .D(D[18]), .CK(net18798), .RN(RST), .Q(Q[18]) );
  DFFR_X1 \Q_reg[17]  ( .D(D[17]), .CK(net18798), .RN(RST), .Q(Q[17]) );
  DFFR_X1 \Q_reg[16]  ( .D(D[16]), .CK(net18798), .RN(RST), .Q(Q[16]) );
  DFFR_X1 \Q_reg[15]  ( .D(D[15]), .CK(net18798), .RN(RST), .Q(Q[15]) );
  DFFR_X1 \Q_reg[14]  ( .D(D[14]), .CK(net18798), .RN(RST), .Q(Q[14]) );
  DFFR_X1 \Q_reg[13]  ( .D(D[13]), .CK(net18798), .RN(RST), .Q(Q[13]) );
  DFFR_X1 \Q_reg[12]  ( .D(D[12]), .CK(net18798), .RN(RST), .Q(Q[12]) );
  DFFR_X1 \Q_reg[11]  ( .D(D[11]), .CK(net18798), .RN(RST), .Q(Q[11]) );
  DFFR_X1 \Q_reg[10]  ( .D(D[10]), .CK(net18798), .RN(RST), .Q(Q[10]) );
  DFFR_X1 \Q_reg[9]  ( .D(D[9]), .CK(net18798), .RN(RST), .Q(Q[9]) );
  DFFR_X1 \Q_reg[8]  ( .D(D[8]), .CK(net18798), .RN(RST), .Q(Q[8]) );
  DFFR_X1 \Q_reg[7]  ( .D(D[7]), .CK(net18798), .RN(RST), .Q(Q[7]) );
  DFFR_X1 \Q_reg[6]  ( .D(D[6]), .CK(net18798), .RN(RST), .Q(Q[6]) );
  DFFR_X1 \Q_reg[5]  ( .D(D[5]), .CK(net18798), .RN(RST), .Q(Q[5]) );
  DFFR_X1 \Q_reg[4]  ( .D(D[4]), .CK(net18798), .RN(RST), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(D[3]), .CK(net18798), .RN(RST), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(n1), .CK(net18798), .RN(RST), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(D[1]), .CK(net18798), .RN(RST), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(D[0]), .CK(net18798), .RN(RST), .Q(Q[0]) );
  INV_X1 U2 ( .A(D[2]), .ZN(n1) );
endmodule


module SNPS_CLOCK_GATE_HIGH_reg_N32_11 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18782, net18784, net18786, net18787, net18790, net18793;
  assign net18782 = EN;
  assign net18784 = CLK;
  assign ENCLK = net18786;
  assign net18793 = TE;

  DLL_X1 latch ( .D(net18787), .GN(net18784), .Q(net18790) );
  AND2_X1 main_gate ( .A1(net18790), .A2(net18784), .ZN(net18786) );
  OR2_X1 test_or ( .A1(net18782), .A2(net18793), .ZN(net18787) );
endmodule


module reg_N32_11 ( D, Q, EN, CLK, RST );
  input [31:0] D;
  output [31:0] Q;
  input EN, CLK, RST;
  wire   net18798;

  SNPS_CLOCK_GATE_HIGH_reg_N32_11 clk_gate_Q_reg ( .CLK(CLK), .EN(EN), .ENCLK(
        net18798), .TE(1'b0) );
  DFFR_X1 \Q_reg[25]  ( .D(D[25]), .CK(net18798), .RN(RST), .Q(Q[25]) );
  DFFR_X1 \Q_reg[24]  ( .D(D[24]), .CK(net18798), .RN(RST), .Q(Q[24]) );
  DFFR_X1 \Q_reg[23]  ( .D(D[23]), .CK(net18798), .RN(RST), .Q(Q[23]) );
  DFFR_X1 \Q_reg[22]  ( .D(D[22]), .CK(net18798), .RN(RST), .Q(Q[22]) );
  DFFR_X1 \Q_reg[21]  ( .D(D[21]), .CK(net18798), .RN(RST), .Q(Q[21]) );
  DFFR_X1 \Q_reg[20]  ( .D(D[20]), .CK(net18798), .RN(RST), .Q(Q[20]) );
  DFFR_X1 \Q_reg[19]  ( .D(D[19]), .CK(net18798), .RN(RST), .Q(Q[19]) );
  DFFR_X1 \Q_reg[18]  ( .D(D[18]), .CK(net18798), .RN(RST), .Q(Q[18]) );
  DFFR_X1 \Q_reg[17]  ( .D(D[17]), .CK(net18798), .RN(RST), .Q(Q[17]) );
  DFFR_X1 \Q_reg[16]  ( .D(D[16]), .CK(net18798), .RN(RST), .Q(Q[16]) );
  DFFR_X1 \Q_reg[15]  ( .D(D[15]), .CK(net18798), .RN(RST), .Q(Q[15]) );
  DFFR_X1 \Q_reg[14]  ( .D(D[14]), .CK(net18798), .RN(RST), .Q(Q[14]) );
  DFFR_X1 \Q_reg[13]  ( .D(D[13]), .CK(net18798), .RN(RST), .Q(Q[13]) );
  DFFR_X1 \Q_reg[12]  ( .D(D[12]), .CK(net18798), .RN(RST), .Q(Q[12]) );
  DFFR_X1 \Q_reg[11]  ( .D(D[11]), .CK(net18798), .RN(RST), .Q(Q[11]) );
  DFFR_X1 \Q_reg[10]  ( .D(D[10]), .CK(net18798), .RN(RST), .Q(Q[10]) );
  DFFR_X1 \Q_reg[9]  ( .D(D[9]), .CK(net18798), .RN(RST), .Q(Q[9]) );
  DFFR_X1 \Q_reg[8]  ( .D(D[8]), .CK(net18798), .RN(RST), .Q(Q[8]) );
  DFFR_X1 \Q_reg[7]  ( .D(D[7]), .CK(net18798), .RN(RST), .Q(Q[7]) );
  DFFR_X1 \Q_reg[6]  ( .D(D[6]), .CK(net18798), .RN(RST), .Q(Q[6]) );
  DFFR_X1 \Q_reg[5]  ( .D(D[5]), .CK(net18798), .RN(RST), .Q(Q[5]) );
  DFFR_X1 \Q_reg[4]  ( .D(D[4]), .CK(net18798), .RN(RST), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(D[3]), .CK(net18798), .RN(RST), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(D[2]), .CK(net18798), .RN(RST), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(D[1]), .CK(net18798), .RN(RST), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(D[0]), .CK(net18798), .RN(RST), .Q(Q[0]) );
endmodule


module MUX_2to1_N32_0 ( IN0, IN1, SEL, Y );
  input [31:0] IN0;
  input [31:0] IN1;
  output [31:0] Y;
  input SEL;
  wire   n1, n2;

  BUF_X1 U1 ( .A(SEL), .Z(n2) );
  BUF_X1 U2 ( .A(SEL), .Z(n1) );
  MUX2_X1 U3 ( .A(IN0[0]), .B(IN1[0]), .S(n1), .Z(Y[0]) );
  MUX2_X1 U4 ( .A(IN0[10]), .B(IN1[10]), .S(n1), .Z(Y[10]) );
  MUX2_X1 U5 ( .A(IN0[11]), .B(IN1[11]), .S(n1), .Z(Y[11]) );
  MUX2_X1 U6 ( .A(IN0[12]), .B(IN1[12]), .S(n1), .Z(Y[12]) );
  MUX2_X1 U7 ( .A(IN0[13]), .B(IN1[13]), .S(n1), .Z(Y[13]) );
  MUX2_X1 U8 ( .A(IN0[14]), .B(IN1[14]), .S(n1), .Z(Y[14]) );
  MUX2_X1 U9 ( .A(IN0[15]), .B(IN1[15]), .S(n1), .Z(Y[15]) );
  MUX2_X1 U10 ( .A(IN0[16]), .B(IN1[16]), .S(n1), .Z(Y[16]) );
  MUX2_X1 U11 ( .A(IN0[17]), .B(IN1[17]), .S(n1), .Z(Y[17]) );
  MUX2_X1 U12 ( .A(IN0[18]), .B(IN1[18]), .S(n1), .Z(Y[18]) );
  MUX2_X1 U13 ( .A(IN0[19]), .B(IN1[19]), .S(n1), .Z(Y[19]) );
  MUX2_X1 U14 ( .A(IN0[1]), .B(IN1[1]), .S(n2), .Z(Y[1]) );
  MUX2_X1 U15 ( .A(IN0[20]), .B(IN1[20]), .S(n2), .Z(Y[20]) );
  MUX2_X1 U16 ( .A(IN0[21]), .B(IN1[21]), .S(n2), .Z(Y[21]) );
  MUX2_X1 U17 ( .A(IN0[22]), .B(IN1[22]), .S(n2), .Z(Y[22]) );
  MUX2_X1 U18 ( .A(IN0[23]), .B(IN1[23]), .S(n2), .Z(Y[23]) );
  MUX2_X1 U19 ( .A(IN0[24]), .B(IN1[24]), .S(n2), .Z(Y[24]) );
  MUX2_X1 U20 ( .A(IN0[25]), .B(IN1[25]), .S(n2), .Z(Y[25]) );
  MUX2_X1 U21 ( .A(IN0[26]), .B(IN1[26]), .S(n2), .Z(Y[26]) );
  MUX2_X1 U22 ( .A(IN0[27]), .B(IN1[27]), .S(n2), .Z(Y[27]) );
  MUX2_X1 U23 ( .A(IN0[28]), .B(IN1[28]), .S(n2), .Z(Y[28]) );
  MUX2_X1 U24 ( .A(IN0[29]), .B(IN1[29]), .S(n2), .Z(Y[29]) );
  MUX2_X1 U25 ( .A(IN0[2]), .B(IN1[2]), .S(n1), .Z(Y[2]) );
  MUX2_X1 U26 ( .A(IN0[30]), .B(IN1[30]), .S(n2), .Z(Y[30]) );
  MUX2_X1 U27 ( .A(IN0[31]), .B(IN1[31]), .S(SEL), .Z(Y[31]) );
  MUX2_X1 U28 ( .A(IN0[3]), .B(IN1[3]), .S(n1), .Z(Y[3]) );
  MUX2_X1 U29 ( .A(IN0[4]), .B(IN1[4]), .S(n2), .Z(Y[4]) );
  MUX2_X1 U30 ( .A(IN0[5]), .B(IN1[5]), .S(SEL), .Z(Y[5]) );
  MUX2_X1 U31 ( .A(IN0[6]), .B(IN1[6]), .S(n1), .Z(Y[6]) );
  MUX2_X1 U32 ( .A(IN0[7]), .B(IN1[7]), .S(SEL), .Z(Y[7]) );
  MUX2_X1 U33 ( .A(IN0[8]), .B(IN1[8]), .S(n1), .Z(Y[8]) );
  MUX2_X1 U34 ( .A(IN0[9]), .B(IN1[9]), .S(n2), .Z(Y[9]) );
endmodule


module PG_NETWORK_0 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_1023 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_1022 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_1021 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_1020 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_1019 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_1018 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_1017 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_1016 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_1015 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_1014 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_1013 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_1012 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_1011 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_1010 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_1009 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_1008 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_1007 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_1006 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_1005 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_1004 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_1003 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_1002 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_1001 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_1000 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_999 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_998 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_997 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module G_BLOCK_0 ( P_ik, G_ik, G_k1j, G_ij );
  input P_ik, G_ik, G_k1j;
  output G_ij;
  wire   n1;

  AOI21_X1 U1 ( .B1(P_ik), .B2(G_k1j), .A(G_ik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_0 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_998 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_997 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_996 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_995 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_994 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_993 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_992 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_991 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_990 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_989 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_988 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_987 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module G_BLOCK_272 ( P_ik, G_ik, G_k1j, G_ij );
  input P_ik, G_ik, G_k1j;
  output G_ij;
  wire   n1;

  AOI21_X1 U1 ( .B1(P_ik), .B2(G_k1j), .A(G_ik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_984 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_983 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_982 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_981 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_980 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_979 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module G_BLOCK_271 ( P_ik, G_ik, G_k1j, G_ij );
  input P_ik, G_ik, G_k1j;
  output G_ij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(G_ij) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(G_k1j), .A(G_ik), .ZN(n1) );
endmodule


module PG_BLOCK_977 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_976 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module G_BLOCK_270 ( P_ik, G_ik, G_k1j, G_ij );
  input P_ik, G_ik, G_k1j;
  output G_ij;
  wire   n1;

  AOI21_X1 U1 ( .B1(P_ik), .B2(G_k1j), .A(G_ik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(G_ij) );
endmodule


module G_BLOCK_269 ( P_ik, G_ik, G_k1j, G_ij );
  input P_ik, G_ik, G_k1j;
  output G_ij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(G_ij) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(G_k1j), .A(G_ik), .ZN(n1) );
endmodule


module PG_BLOCK_974 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module G_BLOCK_268 ( P_ik, G_ik, G_k1j, G_ij );
  input P_ik, G_ik, G_k1j;
  output G_ij;
  wire   n1;

  AOI21_X1 U1 ( .B1(P_ik), .B2(G_k1j), .A(G_ik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(G_ij) );
endmodule


module G_BLOCK_267 ( P_ik, G_ik, G_k1j, G_ij );
  input P_ik, G_ik, G_k1j;
  output G_ij;
  wire   n1;

  AOI21_X1 U1 ( .B1(P_ik), .B2(G_k1j), .A(G_ik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(G_ij) );
endmodule


module G_BLOCK_266 ( P_ik, G_ik, G_k1j, G_ij );
  input P_ik, G_ik, G_k1j;
  output G_ij;
  wire   n1;

  AOI21_X1 U1 ( .B1(P_ik), .B2(G_k1j), .A(G_ik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(G_ij) );
endmodule


module CARRY_GENERATOR_Nbit32_0 ( A, B, Cin, Cout );
  input [31:0] A;
  input [31:0] B;
  output [8:0] Cout;
  input Cin;
  wire   \p[4][2] , \p[3][2] , \p[3][1] , \p[2][6] , \p[2][5] , \p[2][4] ,
         \p[2][3] , \p[2][2] , \p[2][1] , \p[1][13] , \p[1][12] , \p[1][11] ,
         \p[1][10] , \p[1][9] , \p[1][8] , \p[1][7] , \p[1][6] , \p[1][5] ,
         \p[1][4] , \p[1][3] , \p[1][2] , \p[1][1] , \p[0][28] , \p[0][27] ,
         \p[0][26] , \p[0][25] , \p[0][24] , \p[0][23] , \p[0][22] ,
         \p[0][21] , \p[0][20] , \p[0][19] , \p[0][18] , \p[0][17] ,
         \p[0][16] , \p[0][15] , \p[0][14] , \p[0][13] , \p[0][12] ,
         \p[0][11] , \p[0][10] , \p[0][9] , \p[0][8] , \p[0][7] , \p[0][6] ,
         \p[0][5] , \p[0][4] , \p[0][3] , \p[0][2] , \g[4][2] , \g[3][2] ,
         \g[3][1] , \g[2][6] , \g[2][5] , \g[2][4] , \g[2][3] , \g[2][2] ,
         \g[2][1] , \g[1][13] , \g[1][12] , \g[1][11] , \g[1][10] , \g[1][9] ,
         \g[1][8] , \g[1][7] , \g[1][6] , \g[1][5] , \g[1][4] , \g[1][3] ,
         \g[1][2] , \g[1][1] , \g[1][0] , \g[0][28] , \g[0][27] , \g[0][26] ,
         \g[0][25] , \g[0][24] , \g[0][23] , \g[0][22] , \g[0][21] ,
         \g[0][20] , \g[0][19] , \g[0][18] , \g[0][17] , \g[0][16] ,
         \g[0][15] , \g[0][14] , \g[0][13] , \g[0][12] , \g[0][11] ,
         \g[0][10] , \g[0][9] , \g[0][8] , \g[0][7] , \g[0][6] , \g[0][5] ,
         \g[0][4] , \g[0][3] , \g[0][2] , \g[0][1] ;

  PG_NETWORK_0 Block_PG_NET_1 ( .op1(A[0]), .op2(B[0]), .g(\g[0][1] ) );
  PG_NETWORK_1023 Block_PG_NET_2 ( .op1(A[1]), .op2(B[1]), .g(\g[0][2] ), .p(
        \p[0][2] ) );
  PG_NETWORK_1022 Block_PG_NET_3 ( .op1(A[2]), .op2(B[2]), .g(\g[0][3] ), .p(
        \p[0][3] ) );
  PG_NETWORK_1021 Block_PG_NET_4 ( .op1(A[3]), .op2(B[3]), .g(\g[0][4] ), .p(
        \p[0][4] ) );
  PG_NETWORK_1020 Block_PG_NET_5 ( .op1(A[4]), .op2(B[4]), .g(\g[0][5] ), .p(
        \p[0][5] ) );
  PG_NETWORK_1019 Block_PG_NET_6 ( .op1(A[5]), .op2(B[5]), .g(\g[0][6] ), .p(
        \p[0][6] ) );
  PG_NETWORK_1018 Block_PG_NET_7 ( .op1(A[6]), .op2(B[6]), .g(\g[0][7] ), .p(
        \p[0][7] ) );
  PG_NETWORK_1017 Block_PG_NET_8 ( .op1(A[7]), .op2(B[7]), .g(\g[0][8] ), .p(
        \p[0][8] ) );
  PG_NETWORK_1016 Block_PG_NET_9 ( .op1(A[8]), .op2(B[8]), .g(\g[0][9] ), .p(
        \p[0][9] ) );
  PG_NETWORK_1015 Block_PG_NET_10 ( .op1(A[9]), .op2(B[9]), .g(\g[0][10] ), 
        .p(\p[0][10] ) );
  PG_NETWORK_1014 Block_PG_NET_11 ( .op1(A[10]), .op2(B[10]), .g(\g[0][11] ), 
        .p(\p[0][11] ) );
  PG_NETWORK_1013 Block_PG_NET_12 ( .op1(A[11]), .op2(B[11]), .g(\g[0][12] ), 
        .p(\p[0][12] ) );
  PG_NETWORK_1012 Block_PG_NET_13 ( .op1(A[12]), .op2(B[12]), .g(\g[0][13] ), 
        .p(\p[0][13] ) );
  PG_NETWORK_1011 Block_PG_NET_14 ( .op1(A[13]), .op2(B[13]), .g(\g[0][14] ), 
        .p(\p[0][14] ) );
  PG_NETWORK_1010 Block_PG_NET_15 ( .op1(A[14]), .op2(B[14]), .g(\g[0][15] ), 
        .p(\p[0][15] ) );
  PG_NETWORK_1009 Block_PG_NET_16 ( .op1(A[15]), .op2(B[15]), .g(\g[0][16] ), 
        .p(\p[0][16] ) );
  PG_NETWORK_1008 Block_PG_NET_17 ( .op1(A[16]), .op2(B[16]), .g(\g[0][17] ), 
        .p(\p[0][17] ) );
  PG_NETWORK_1007 Block_PG_NET_18 ( .op1(A[17]), .op2(B[17]), .g(\g[0][18] ), 
        .p(\p[0][18] ) );
  PG_NETWORK_1006 Block_PG_NET_19 ( .op1(A[18]), .op2(B[18]), .g(\g[0][19] ), 
        .p(\p[0][19] ) );
  PG_NETWORK_1005 Block_PG_NET_20 ( .op1(A[19]), .op2(B[19]), .g(\g[0][20] ), 
        .p(\p[0][20] ) );
  PG_NETWORK_1004 Block_PG_NET_21 ( .op1(A[20]), .op2(B[20]), .g(\g[0][21] ), 
        .p(\p[0][21] ) );
  PG_NETWORK_1003 Block_PG_NET_22 ( .op1(A[21]), .op2(B[21]), .g(\g[0][22] ), 
        .p(\p[0][22] ) );
  PG_NETWORK_1002 Block_PG_NET_23 ( .op1(A[22]), .op2(B[22]), .g(\g[0][23] ), 
        .p(\p[0][23] ) );
  PG_NETWORK_1001 Block_PG_NET_24 ( .op1(A[23]), .op2(B[23]), .g(\g[0][24] ), 
        .p(\p[0][24] ) );
  PG_NETWORK_1000 Block_PG_NET_25 ( .op1(A[24]), .op2(B[24]), .g(\g[0][25] ), 
        .p(\p[0][25] ) );
  PG_NETWORK_999 Block_PG_NET_26 ( .op1(A[25]), .op2(B[25]), .g(\g[0][26] ), 
        .p(\p[0][26] ) );
  PG_NETWORK_998 Block_PG_NET_27 ( .op1(A[26]), .op2(B[26]), .g(\g[0][27] ), 
        .p(\p[0][27] ) );
  PG_NETWORK_997 Block_PG_NET_28 ( .op1(A[27]), .op2(B[27]), .g(\g[0][28] ), 
        .p(\p[0][28] ) );
  G_BLOCK_0 g_1 ( .P_ik(\p[0][2] ), .G_ik(\g[0][2] ), .G_k1j(\g[0][1] ), 
        .G_ij(\g[1][0] ) );
  PG_BLOCK_0 Block_Stage_ONE_1 ( .P_ik(\p[0][4] ), .G_ik(\g[0][4] ), .P_k1j(
        \p[0][3] ), .G_k1j(\g[0][3] ), .P_ij(\p[1][1] ), .G_ij(\g[1][1] ) );
  PG_BLOCK_998 Block_Stage_ONE_2 ( .P_ik(\p[0][6] ), .G_ik(\g[0][6] ), .P_k1j(
        \p[0][5] ), .G_k1j(\g[0][5] ), .P_ij(\p[1][2] ), .G_ij(\g[1][2] ) );
  PG_BLOCK_997 Block_Stage_ONE_3 ( .P_ik(\p[0][8] ), .G_ik(\g[0][8] ), .P_k1j(
        \p[0][7] ), .G_k1j(\g[0][7] ), .P_ij(\p[1][3] ), .G_ij(\g[1][3] ) );
  PG_BLOCK_996 Block_Stage_ONE_4 ( .P_ik(\p[0][10] ), .G_ik(\g[0][10] ), 
        .P_k1j(\p[0][9] ), .G_k1j(\g[0][9] ), .P_ij(\p[1][4] ), .G_ij(
        \g[1][4] ) );
  PG_BLOCK_995 Block_Stage_ONE_5 ( .P_ik(\p[0][12] ), .G_ik(\g[0][12] ), 
        .P_k1j(\p[0][11] ), .G_k1j(\g[0][11] ), .P_ij(\p[1][5] ), .G_ij(
        \g[1][5] ) );
  PG_BLOCK_994 Block_Stage_ONE_6 ( .P_ik(\p[0][14] ), .G_ik(\g[0][14] ), 
        .P_k1j(\p[0][13] ), .G_k1j(\g[0][13] ), .P_ij(\p[1][6] ), .G_ij(
        \g[1][6] ) );
  PG_BLOCK_993 Block_Stage_ONE_7 ( .P_ik(\p[0][16] ), .G_ik(\g[0][16] ), 
        .P_k1j(\p[0][15] ), .G_k1j(\g[0][15] ), .P_ij(\p[1][7] ), .G_ij(
        \g[1][7] ) );
  PG_BLOCK_992 Block_Stage_ONE_8 ( .P_ik(\p[0][18] ), .G_ik(\g[0][18] ), 
        .P_k1j(\p[0][17] ), .G_k1j(\g[0][17] ), .P_ij(\p[1][8] ), .G_ij(
        \g[1][8] ) );
  PG_BLOCK_991 Block_Stage_ONE_9 ( .P_ik(\p[0][20] ), .G_ik(\g[0][20] ), 
        .P_k1j(\p[0][19] ), .G_k1j(\g[0][19] ), .P_ij(\p[1][9] ), .G_ij(
        \g[1][9] ) );
  PG_BLOCK_990 Block_Stage_ONE_10 ( .P_ik(\p[0][22] ), .G_ik(\g[0][22] ), 
        .P_k1j(\p[0][21] ), .G_k1j(\g[0][21] ), .P_ij(\p[1][10] ), .G_ij(
        \g[1][10] ) );
  PG_BLOCK_989 Block_Stage_ONE_11 ( .P_ik(\p[0][24] ), .G_ik(\g[0][24] ), 
        .P_k1j(\p[0][23] ), .G_k1j(\g[0][23] ), .P_ij(\p[1][11] ), .G_ij(
        \g[1][11] ) );
  PG_BLOCK_988 Block_Stage_ONE_12 ( .P_ik(\p[0][26] ), .G_ik(\g[0][26] ), 
        .P_k1j(\p[0][25] ), .G_k1j(\g[0][25] ), .P_ij(\p[1][12] ), .G_ij(
        \g[1][12] ) );
  PG_BLOCK_987 Block_Stage_ONE_13 ( .P_ik(\p[0][28] ), .G_ik(\g[0][28] ), 
        .P_k1j(\p[0][27] ), .G_k1j(\g[0][27] ), .P_ij(\p[1][13] ), .G_ij(
        \g[1][13] ) );
  G_BLOCK_272 g_2 ( .P_ik(\p[1][1] ), .G_ik(\g[1][1] ), .G_k1j(\g[1][0] ), 
        .G_ij(Cout[1]) );
  PG_BLOCK_984 Block_Stage_TWO_1 ( .P_ik(\p[1][3] ), .G_ik(\g[1][3] ), .P_k1j(
        \p[1][2] ), .G_k1j(\g[1][2] ), .P_ij(\p[2][1] ), .G_ij(\g[2][1] ) );
  PG_BLOCK_983 Block_Stage_TWO_2 ( .P_ik(\p[1][5] ), .G_ik(\g[1][5] ), .P_k1j(
        \p[1][4] ), .G_k1j(\g[1][4] ), .P_ij(\p[2][2] ), .G_ij(\g[2][2] ) );
  PG_BLOCK_982 Block_Stage_TWO_3 ( .P_ik(\p[1][7] ), .G_ik(\g[1][7] ), .P_k1j(
        \p[1][6] ), .G_k1j(\g[1][6] ), .P_ij(\p[2][3] ), .G_ij(\g[2][3] ) );
  PG_BLOCK_981 Block_Stage_TWO_4 ( .P_ik(\p[1][9] ), .G_ik(\g[1][9] ), .P_k1j(
        \p[1][8] ), .G_k1j(\g[1][8] ), .P_ij(\p[2][4] ), .G_ij(\g[2][4] ) );
  PG_BLOCK_980 Block_Stage_TWO_5 ( .P_ik(\p[1][11] ), .G_ik(\g[1][11] ), 
        .P_k1j(\p[1][10] ), .G_k1j(\g[1][10] ), .P_ij(\p[2][5] ), .G_ij(
        \g[2][5] ) );
  PG_BLOCK_979 Block_Stage_TWO_6 ( .P_ik(\p[1][13] ), .G_ik(\g[1][13] ), 
        .P_k1j(\p[1][12] ), .G_k1j(\g[1][12] ), .P_ij(\p[2][6] ), .G_ij(
        \g[2][6] ) );
  G_BLOCK_271 g_3 ( .P_ik(\p[2][1] ), .G_ik(\g[2][1] ), .G_k1j(Cout[1]), 
        .G_ij(Cout[2]) );
  PG_BLOCK_977 Block_Stage_THREE_1 ( .P_ik(\p[2][3] ), .G_ik(\g[2][3] ), 
        .P_k1j(\p[2][2] ), .G_k1j(\g[2][2] ), .P_ij(\p[3][1] ), .G_ij(
        \g[3][1] ) );
  PG_BLOCK_976 Block_Stage_THREE_2 ( .P_ik(\p[2][5] ), .G_ik(\g[2][5] ), 
        .P_k1j(\p[2][4] ), .G_k1j(\g[2][4] ), .P_ij(\p[3][2] ), .G_ij(
        \g[3][2] ) );
  G_BLOCK_270 g_4_c12_c16_0 ( .P_ik(\p[2][2] ), .G_ik(\g[2][2] ), .G_k1j(
        Cout[2]), .G_ij(Cout[3]) );
  G_BLOCK_269 g_4_c12_c16_1 ( .P_ik(\p[3][1] ), .G_ik(\g[3][1] ), .G_k1j(
        Cout[2]), .G_ij(Cout[4]) );
  PG_BLOCK_974 Block_stage_FOUR_2_0 ( .P_ik(\p[2][6] ), .G_ik(\g[2][6] ), 
        .P_k1j(\p[3][2] ), .G_k1j(\g[3][2] ), .P_ij(\p[4][2] ), .G_ij(
        \g[4][2] ) );
  G_BLOCK_268 Block_stage_FIVE_4 ( .P_ik(\p[2][4] ), .G_ik(\g[2][4] ), .G_k1j(
        Cout[4]), .G_ij(Cout[5]) );
  G_BLOCK_267 Block_stage_FIVE_5 ( .P_ik(\p[3][2] ), .G_ik(\g[3][2] ), .G_k1j(
        Cout[4]), .G_ij(Cout[6]) );
  G_BLOCK_266 Block_stage_FIVE_6 ( .P_ik(\p[4][2] ), .G_ik(\g[4][2] ), .G_k1j(
        Cout[4]), .G_ij(Cout[7]) );
endmodule


module FA_2048 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_2047 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_2046 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_2045 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_0 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_2048 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_2047 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_2046 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_2045 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_256 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_0 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_0 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  MUX_2to1_N4_256 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_2040 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_2039 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_2038 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_2037 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_510 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_2040 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_2039 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_2038 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_2037 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_2036 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_2035 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_2034 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_2033 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_509 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_2036 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_2035 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_2034 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_2033 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_255 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U3 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U4 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
endmodule


module carry_select_block_N4_255 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_510 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_509 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_255 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_2032 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_2031 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_2030 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_2029 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_508 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_2032 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_2031 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_2030 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_2029 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_2028 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_2027 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_2026 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_2025 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_507 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_2028 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_2027 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_2026 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_2025 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_254 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U3 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U4 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
endmodule


module carry_select_block_N4_254 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_508 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_507 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_254 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_2024 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_2023 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_2022 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_2021 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_506 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_2024 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_2023 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_2022 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_2021 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_2020 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_2019 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_2018 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_2017 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_505 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_2020 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_2019 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_2018 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_2017 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_253 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U3 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U4 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
endmodule


module carry_select_block_N4_253 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_506 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_505 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_253 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_2016 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_2015 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_2014 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_2013 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_504 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_2016 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_2015 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_2014 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_2013 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_2012 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_2011 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_2010 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_2009 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_503 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_2012 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_2011 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_2010 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_2009 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_252 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U3 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U4 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
endmodule


module carry_select_block_N4_252 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_504 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_503 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_252 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_2008 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_2007 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_2006 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_2005 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_502 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_2008 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_2007 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_2006 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_2005 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_2004 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_2003 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_2002 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_2001 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_501 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_2004 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_2003 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_2002 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_2001 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_251 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U3 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U4 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
endmodule


module carry_select_block_N4_251 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_502 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_501 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_251 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_2000 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1999 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1998 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1997 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n2) );
  XNOR2_X1 U2 ( .A(n2), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_500 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_2000 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1999 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1998 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1997 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1996 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_1995 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1994 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1993 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n2) );
  XNOR2_X1 U2 ( .A(n2), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_499 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1996 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1995 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1994 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1993 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_250 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U3 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U4 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
endmodule


module carry_select_block_N4_250 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_500 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_499 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_250 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_1992 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1991 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1990 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1989 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n2) );
  XNOR2_X1 U2 ( .A(n2), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_498 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1992 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1991 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1990 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1989 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1988 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_1987 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1986 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1985 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n2) );
  XNOR2_X1 U2 ( .A(n2), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_497 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1988 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1987 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1986 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1985 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_249 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U3 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U4 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
endmodule


module carry_select_block_N4_249 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_498 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_497 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_249 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module SUMGENERATOR_Nblocks8_bits_per_block4_0 ( A, B, CARRY_SELECT, SUM );
  input [31:0] A;
  input [31:0] B;
  input [7:0] CARRY_SELECT;
  output [31:0] SUM;


  carry_select_block_N4_0 block_n_1 ( .A(A[3:0]), .B(B[3:0]), .S(SUM[3:0]), 
        .Ci(1'b0) );
  carry_select_block_N4_255 block_n_2 ( .A(A[7:4]), .B(B[7:4]), .S(SUM[7:4]), 
        .Ci(CARRY_SELECT[1]) );
  carry_select_block_N4_254 block_n_3 ( .A(A[11:8]), .B(B[11:8]), .S(SUM[11:8]), .Ci(CARRY_SELECT[2]) );
  carry_select_block_N4_253 block_n_4 ( .A(A[15:12]), .B(B[15:12]), .S(
        SUM[15:12]), .Ci(CARRY_SELECT[3]) );
  carry_select_block_N4_252 block_n_5 ( .A(A[19:16]), .B(B[19:16]), .S(
        SUM[19:16]), .Ci(CARRY_SELECT[4]) );
  carry_select_block_N4_251 block_n_6 ( .A(A[23:20]), .B(B[23:20]), .S(
        SUM[23:20]), .Ci(CARRY_SELECT[5]) );
  carry_select_block_N4_250 block_n_7 ( .A(A[27:24]), .B(B[27:24]), .S(
        SUM[27:24]), .Ci(CARRY_SELECT[6]) );
  carry_select_block_N4_249 block_n_8 ( .A(A[31:28]), .B(B[31:28]), .S(
        SUM[31:28]), .Ci(CARRY_SELECT[7]) );
endmodule


module ADDER_P4_N_BIT32_0 ( A, B, add_sub, Cout, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input add_sub;
  output Cout;

  wire   [31:0] B_xor;
  wire   [7:0] tmp_co;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign B_xor[24] = B[24];
  assign B_xor[23] = B[23];
  assign B_xor[22] = B[22];
  assign B_xor[21] = B[21];
  assign B_xor[20] = B[20];
  assign B_xor[19] = B[19];
  assign B_xor[18] = B[18];
  assign B_xor[17] = B[17];
  assign B_xor[16] = B[16];
  assign B_xor[15] = B[15];
  assign B_xor[14] = B[14];
  assign B_xor[13] = B[13];
  assign B_xor[12] = B[12];
  assign B_xor[11] = B[11];
  assign B_xor[10] = B[10];
  assign B_xor[9] = B[9];
  assign B_xor[8] = B[8];
  assign B_xor[7] = B[7];
  assign B_xor[6] = B[6];
  assign B_xor[5] = B[5];
  assign B_xor[4] = B[4];
  assign B_xor[3] = B[3];
  assign B_xor[2] = B[2];
  assign B_xor[1] = B[1];
  assign B_xor[0] = B[0];

  CARRY_GENERATOR_Nbit32_0 CLA_SPARSE_TREE ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        A[27:0]}), .B({1'b0, 1'b0, 1'b0, 1'b0, B[27:25], B_xor[24:0]}), .Cin(
        1'b0), .Cout({SYNOPSYS_UNCONNECTED__0, tmp_co[7:1], 
        SYNOPSYS_UNCONNECTED__1}) );
  SUMGENERATOR_Nblocks8_bits_per_block4_0 CSA ( .A(A), .B({B[31:25], 
        B_xor[24:0]}), .CARRY_SELECT({tmp_co[7:1], 1'b0}), .SUM(SUM) );
endmodule


module branch_comp_N32 ( .BRANCH_COND({\BRANCH_COND[1] , \BRANCH_COND[0] }), 
        DATA_IN, BRANCH_IS_TAKEN );
  input [31:0] DATA_IN;
  input \BRANCH_COND[1] , \BRANCH_COND[0] ;
  output BRANCH_IS_TAKEN;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19;
  wire   [1:0] BRANCH_COND;

  NAND3_X1 U3 ( .A1(n2), .A2(n1), .A3(n3), .ZN(n7) );
  AND3_X1 U4 ( .A1(n14), .A2(n15), .A3(BRANCH_COND[1]), .ZN(n1) );
  AND4_X1 U5 ( .A1(n19), .A2(n18), .A3(n16), .A4(n10), .ZN(n2) );
  NOR4_X1 U6 ( .A1(DATA_IN[30]), .A2(DATA_IN[3]), .A3(DATA_IN[13]), .A4(
        DATA_IN[14]), .ZN(n3) );
  INV_X1 U7 ( .A(DATA_IN[7]), .ZN(n4) );
  INV_X1 U8 ( .A(DATA_IN[9]), .ZN(n5) );
  INV_X1 U9 ( .A(DATA_IN[10]), .ZN(n6) );
  NAND3_X1 U10 ( .A1(n6), .A2(n5), .A3(n4), .ZN(n13) );
  XNOR2_X1 U11 ( .A(n8), .B(n9), .ZN(BRANCH_IS_TAKEN) );
  NOR2_X1 U12 ( .A1(n7), .A2(DATA_IN[0]), .ZN(n8) );
  INV_X1 U13 ( .A(BRANCH_COND[0]), .ZN(n9) );
  AND2_X1 U14 ( .A1(n17), .A2(n11), .ZN(n10) );
  NOR2_X1 U15 ( .A1(n13), .A2(n12), .ZN(n11) );
  OR2_X1 U16 ( .A1(DATA_IN[11]), .A2(DATA_IN[12]), .ZN(n12) );
  NOR4_X1 U17 ( .A1(DATA_IN[4]), .A2(DATA_IN[5]), .A3(DATA_IN[6]), .A4(
        DATA_IN[8]), .ZN(n15) );
  NOR2_X1 U18 ( .A1(DATA_IN[31]), .A2(DATA_IN[2]), .ZN(n14) );
  NOR4_X1 U19 ( .A1(DATA_IN[26]), .A2(DATA_IN[27]), .A3(DATA_IN[28]), .A4(
        DATA_IN[29]), .ZN(n18) );
  NOR4_X1 U20 ( .A1(DATA_IN[15]), .A2(DATA_IN[16]), .A3(DATA_IN[17]), .A4(
        DATA_IN[18]), .ZN(n17) );
  NOR4_X1 U21 ( .A1(DATA_IN[22]), .A2(DATA_IN[23]), .A3(DATA_IN[24]), .A4(
        DATA_IN[25]), .ZN(n16) );
  NOR4_X1 U22 ( .A1(DATA_IN[19]), .A2(DATA_IN[1]), .A3(DATA_IN[20]), .A4(
        DATA_IN[21]), .ZN(n19) );
endmodule


module MUX_2to1_N32_9 ( IN0, IN1, SEL, Y );
  input [31:0] IN0;
  input [31:0] IN1;
  output [31:0] Y;
  input SEL;
  wire   n1, n2, n3, n4, n5;

  MUX2_X1 U1 ( .A(IN0[22]), .B(IN1[22]), .S(n5), .Z(Y[22]) );
  CLKBUF_X3 U2 ( .A(SEL), .Z(n3) );
  BUF_X2 U3 ( .A(SEL), .Z(n4) );
  OAI21_X1 U4 ( .B1(n3), .B2(n2), .A(n1), .ZN(Y[18]) );
  NAND2_X1 U5 ( .A1(n5), .A2(IN1[18]), .ZN(n1) );
  INV_X1 U6 ( .A(IN0[18]), .ZN(n2) );
  CLKBUF_X3 U7 ( .A(SEL), .Z(n5) );
  MUX2_X1 U8 ( .A(IN0[0]), .B(IN1[0]), .S(n5), .Z(Y[0]) );
  MUX2_X1 U9 ( .A(IN0[10]), .B(IN1[10]), .S(n4), .Z(Y[10]) );
  MUX2_X1 U10 ( .A(IN0[11]), .B(IN1[11]), .S(n4), .Z(Y[11]) );
  MUX2_X1 U11 ( .A(IN0[12]), .B(IN1[12]), .S(n3), .Z(Y[12]) );
  MUX2_X1 U12 ( .A(IN0[13]), .B(IN1[13]), .S(n5), .Z(Y[13]) );
  MUX2_X1 U13 ( .A(IN0[14]), .B(IN1[14]), .S(n3), .Z(Y[14]) );
  MUX2_X1 U14 ( .A(IN0[15]), .B(IN1[15]), .S(n5), .Z(Y[15]) );
  MUX2_X1 U15 ( .A(IN0[16]), .B(IN1[16]), .S(n3), .Z(Y[16]) );
  MUX2_X1 U16 ( .A(IN0[17]), .B(IN1[17]), .S(n3), .Z(Y[17]) );
  MUX2_X1 U17 ( .A(IN0[19]), .B(IN1[19]), .S(n5), .Z(Y[19]) );
  MUX2_X1 U18 ( .A(IN0[1]), .B(IN1[1]), .S(n3), .Z(Y[1]) );
  MUX2_X1 U19 ( .A(IN0[20]), .B(IN1[20]), .S(n4), .Z(Y[20]) );
  MUX2_X1 U20 ( .A(IN0[21]), .B(IN1[21]), .S(n3), .Z(Y[21]) );
  MUX2_X1 U21 ( .A(IN0[23]), .B(IN1[23]), .S(n5), .Z(Y[23]) );
  MUX2_X1 U22 ( .A(IN0[24]), .B(IN1[24]), .S(n4), .Z(Y[24]) );
  MUX2_X1 U23 ( .A(IN0[25]), .B(IN1[25]), .S(n5), .Z(Y[25]) );
  MUX2_X1 U24 ( .A(IN0[26]), .B(IN1[26]), .S(n4), .Z(Y[26]) );
  MUX2_X1 U25 ( .A(IN0[27]), .B(IN1[27]), .S(n4), .Z(Y[27]) );
  MUX2_X1 U26 ( .A(IN0[28]), .B(IN1[28]), .S(n4), .Z(Y[28]) );
  MUX2_X1 U27 ( .A(IN0[29]), .B(IN1[29]), .S(n3), .Z(Y[29]) );
  MUX2_X1 U28 ( .A(IN0[2]), .B(IN1[2]), .S(n5), .Z(Y[2]) );
  MUX2_X1 U29 ( .A(IN0[30]), .B(IN1[30]), .S(n3), .Z(Y[30]) );
  MUX2_X1 U30 ( .A(IN0[31]), .B(IN1[31]), .S(n3), .Z(Y[31]) );
  MUX2_X1 U31 ( .A(IN0[3]), .B(IN1[3]), .S(n5), .Z(Y[3]) );
  MUX2_X1 U32 ( .A(IN0[4]), .B(IN1[4]), .S(n4), .Z(Y[4]) );
  MUX2_X1 U33 ( .A(IN0[5]), .B(IN1[5]), .S(n4), .Z(Y[5]) );
  MUX2_X1 U34 ( .A(IN0[6]), .B(IN1[6]), .S(n3), .Z(Y[6]) );
  MUX2_X1 U35 ( .A(IN0[7]), .B(IN1[7]), .S(n4), .Z(Y[7]) );
  MUX2_X1 U36 ( .A(IN0[8]), .B(IN1[8]), .S(n3), .Z(Y[8]) );
  MUX2_X1 U37 ( .A(IN0[9]), .B(IN1[9]), .S(n4), .Z(Y[9]) );
endmodule


module MUX_8to1_N32_0 ( IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, SEL, Y );
  input [31:0] IN0;
  input [31:0] IN1;
  input [31:0] IN2;
  input [31:0] IN3;
  input [31:0] IN4;
  input [31:0] IN5;
  input [31:0] IN6;
  input [31:0] IN7;
  input [2:0] SEL;
  output [31:0] Y;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189;

  AND2_X1 U1 ( .A1(n96), .A2(n94), .ZN(n1) );
  AOI22_X1 U2 ( .A1(n9), .A2(IN1[10]), .B1(IN0[10]), .B2(n61), .ZN(n48) );
  AOI22_X1 U3 ( .A1(IN1[11]), .A2(n9), .B1(IN0[11]), .B2(n61), .ZN(n47) );
  AOI22_X1 U4 ( .A1(n8), .A2(IN2[30]), .B1(n7), .B2(IN3[30]), .ZN(n2) );
  AOI22_X1 U5 ( .A1(n11), .A2(IN4[30]), .B1(n6), .B2(IN6[30]), .ZN(n3) );
  AOI22_X1 U6 ( .A1(n10), .A2(IN0[30]), .B1(n12), .B2(IN5[30]), .ZN(n4) );
  NAND2_X1 U7 ( .A1(n9), .A2(IN1[30]), .ZN(n5) );
  NAND4_X1 U8 ( .A1(n2), .A2(n3), .A3(n4), .A4(n5), .ZN(Y[30]) );
  NAND3_X1 U9 ( .A1(n97), .A2(n95), .A3(n1), .ZN(Y[17]) );
  BUF_X2 U10 ( .A(n185), .Z(n6) );
  BUF_X2 U11 ( .A(n182), .Z(n7) );
  BUF_X2 U12 ( .A(n183), .Z(n8) );
  BUF_X2 U13 ( .A(n180), .Z(n9) );
  BUF_X2 U14 ( .A(n181), .Z(n10) );
  BUF_X2 U15 ( .A(n184), .Z(n11) );
  BUF_X2 U16 ( .A(n186), .Z(n12) );
  BUF_X1 U17 ( .A(n181), .Z(n61) );
  NAND4_X1 U18 ( .A1(n45), .A2(n187), .A3(n188), .A4(n189), .ZN(Y[9]) );
  AOI21_X1 U19 ( .B1(IN1[9]), .B2(n9), .A(n46), .ZN(n45) );
  AND2_X1 U20 ( .A1(n10), .A2(IN0[9]), .ZN(n46) );
  NAND4_X1 U21 ( .A1(n73), .A2(n71), .A3(n72), .A4(n47), .ZN(Y[11]) );
  NAND4_X1 U22 ( .A1(n48), .A2(n68), .A3(n69), .A4(n70), .ZN(Y[10]) );
  NAND4_X1 U23 ( .A1(n175), .A2(n173), .A3(n174), .A4(n49), .ZN(Y[7]) );
  AOI21_X1 U24 ( .B1(n9), .B2(IN1[7]), .A(n50), .ZN(n49) );
  AND2_X1 U25 ( .A1(n10), .A2(IN0[7]), .ZN(n50) );
  NAND2_X1 U26 ( .A1(n55), .A2(n56), .ZN(Y[0]) );
  NOR3_X1 U27 ( .A1(n60), .A2(n59), .A3(n57), .ZN(n56) );
  NAND2_X1 U28 ( .A1(IN1[0]), .A2(n9), .ZN(n55) );
  NOR3_X1 U29 ( .A1(SEL[1]), .A2(n64), .A3(n63), .ZN(n186) );
  INV_X1 U30 ( .A(SEL[2]), .ZN(n63) );
  INV_X1 U31 ( .A(SEL[0]), .ZN(n64) );
  INV_X1 U32 ( .A(SEL[1]), .ZN(n62) );
  INV_X1 U33 ( .A(n51), .ZN(Y[31]) );
  AOI21_X1 U34 ( .B1(IN1[31]), .B2(n9), .A(n52), .ZN(n51) );
  AND2_X1 U35 ( .A1(n154), .A2(n54), .ZN(n53) );
  NAND2_X1 U36 ( .A1(n10), .A2(IN0[31]), .ZN(n54) );
  NAND2_X1 U37 ( .A1(n65), .A2(n58), .ZN(n57) );
  NAND2_X1 U38 ( .A1(n61), .A2(IN0[0]), .ZN(n58) );
  INV_X1 U39 ( .A(n66), .ZN(n59) );
  INV_X1 U40 ( .A(n67), .ZN(n60) );
  NAND3_X1 U41 ( .A1(n156), .A2(n155), .A3(n53), .ZN(n52) );
  NOR3_X1 U42 ( .A1(SEL[2]), .A2(SEL[0]), .A3(SEL[1]), .ZN(n181) );
  NOR3_X1 U43 ( .A1(SEL[2]), .A2(SEL[1]), .A3(n64), .ZN(n180) );
  NOR3_X1 U44 ( .A1(SEL[2]), .A2(SEL[0]), .A3(n62), .ZN(n183) );
  NOR3_X1 U45 ( .A1(SEL[2]), .A2(n64), .A3(n62), .ZN(n182) );
  AOI22_X1 U46 ( .A1(n8), .A2(IN2[0]), .B1(n7), .B2(IN3[0]), .ZN(n67) );
  NOR3_X1 U47 ( .A1(SEL[0]), .A2(n63), .A3(n62), .ZN(n185) );
  NOR3_X1 U48 ( .A1(SEL[0]), .A2(SEL[1]), .A3(n63), .ZN(n184) );
  AOI22_X1 U49 ( .A1(n6), .A2(IN6[0]), .B1(n11), .B2(IN4[0]), .ZN(n66) );
  NAND2_X1 U50 ( .A1(n12), .A2(IN5[0]), .ZN(n65) );
  AOI22_X1 U51 ( .A1(n8), .A2(IN2[10]), .B1(n7), .B2(IN3[10]), .ZN(n70) );
  AOI22_X1 U52 ( .A1(n6), .A2(IN6[10]), .B1(n11), .B2(IN4[10]), .ZN(n69) );
  NAND2_X1 U53 ( .A1(n12), .A2(IN5[10]), .ZN(n68) );
  AOI22_X1 U54 ( .A1(n8), .A2(IN2[11]), .B1(n7), .B2(IN3[11]), .ZN(n73) );
  AOI22_X1 U55 ( .A1(n6), .A2(IN6[11]), .B1(n11), .B2(IN4[11]), .ZN(n72) );
  NAND2_X1 U56 ( .A1(n12), .A2(IN5[11]), .ZN(n71) );
  AOI22_X1 U57 ( .A1(n61), .A2(IN0[12]), .B1(n9), .B2(IN1[12]), .ZN(n77) );
  AOI22_X1 U58 ( .A1(n8), .A2(IN2[12]), .B1(n7), .B2(IN3[12]), .ZN(n76) );
  AOI22_X1 U59 ( .A1(n6), .A2(IN6[12]), .B1(n11), .B2(IN4[12]), .ZN(n75) );
  NAND2_X1 U60 ( .A1(n12), .A2(IN5[12]), .ZN(n74) );
  NAND4_X1 U61 ( .A1(n77), .A2(n76), .A3(n75), .A4(n74), .ZN(Y[12]) );
  AOI22_X1 U62 ( .A1(n61), .A2(IN0[13]), .B1(n9), .B2(IN1[13]), .ZN(n81) );
  AOI22_X1 U63 ( .A1(n8), .A2(IN2[13]), .B1(n7), .B2(IN3[13]), .ZN(n80) );
  AOI22_X1 U64 ( .A1(n6), .A2(IN6[13]), .B1(n11), .B2(IN4[13]), .ZN(n79) );
  NAND2_X1 U65 ( .A1(n12), .A2(IN5[13]), .ZN(n78) );
  NAND4_X1 U66 ( .A1(n81), .A2(n80), .A3(n79), .A4(n78), .ZN(Y[13]) );
  AOI22_X1 U67 ( .A1(n61), .A2(IN0[14]), .B1(n9), .B2(IN1[14]), .ZN(n85) );
  AOI22_X1 U68 ( .A1(n8), .A2(IN2[14]), .B1(n7), .B2(IN3[14]), .ZN(n84) );
  AOI22_X1 U69 ( .A1(n6), .A2(IN6[14]), .B1(n11), .B2(IN4[14]), .ZN(n83) );
  NAND2_X1 U70 ( .A1(n12), .A2(IN5[14]), .ZN(n82) );
  NAND4_X1 U71 ( .A1(n85), .A2(n84), .A3(n83), .A4(n82), .ZN(Y[14]) );
  AOI22_X1 U72 ( .A1(n61), .A2(IN0[15]), .B1(n9), .B2(IN1[15]), .ZN(n89) );
  AOI22_X1 U73 ( .A1(n8), .A2(IN2[15]), .B1(n7), .B2(IN3[15]), .ZN(n88) );
  AOI22_X1 U74 ( .A1(n6), .A2(IN6[15]), .B1(n11), .B2(IN4[15]), .ZN(n87) );
  NAND2_X1 U75 ( .A1(n12), .A2(IN5[15]), .ZN(n86) );
  NAND4_X1 U76 ( .A1(n89), .A2(n88), .A3(n87), .A4(n86), .ZN(Y[15]) );
  AOI22_X1 U77 ( .A1(n61), .A2(IN0[16]), .B1(n9), .B2(IN1[16]), .ZN(n93) );
  AOI22_X1 U78 ( .A1(n8), .A2(IN2[16]), .B1(n7), .B2(IN3[16]), .ZN(n92) );
  AOI22_X1 U79 ( .A1(n6), .A2(IN6[16]), .B1(n11), .B2(IN4[16]), .ZN(n91) );
  NAND2_X1 U80 ( .A1(n12), .A2(IN5[16]), .ZN(n90) );
  NAND4_X1 U81 ( .A1(n93), .A2(n92), .A3(n91), .A4(n90), .ZN(Y[16]) );
  AOI22_X1 U82 ( .A1(n61), .A2(IN0[17]), .B1(n9), .B2(IN1[17]), .ZN(n97) );
  AOI22_X1 U83 ( .A1(n8), .A2(IN2[17]), .B1(n7), .B2(IN3[17]), .ZN(n96) );
  AOI22_X1 U84 ( .A1(n6), .A2(IN6[17]), .B1(n11), .B2(IN4[17]), .ZN(n95) );
  NAND2_X1 U85 ( .A1(n12), .A2(IN5[17]), .ZN(n94) );
  AOI22_X1 U86 ( .A1(n61), .A2(IN0[18]), .B1(n9), .B2(IN1[18]), .ZN(n101) );
  AOI22_X1 U87 ( .A1(n8), .A2(IN2[18]), .B1(n7), .B2(IN3[18]), .ZN(n100) );
  AOI22_X1 U88 ( .A1(n6), .A2(IN6[18]), .B1(n11), .B2(IN4[18]), .ZN(n99) );
  NAND2_X1 U89 ( .A1(n12), .A2(IN5[18]), .ZN(n98) );
  NAND4_X1 U90 ( .A1(n101), .A2(n100), .A3(n99), .A4(n98), .ZN(Y[18]) );
  AOI22_X1 U91 ( .A1(n61), .A2(IN0[19]), .B1(n9), .B2(IN1[19]), .ZN(n105) );
  AOI22_X1 U92 ( .A1(n8), .A2(IN2[19]), .B1(n7), .B2(IN3[19]), .ZN(n104) );
  AOI22_X1 U93 ( .A1(n6), .A2(IN6[19]), .B1(n11), .B2(IN4[19]), .ZN(n103) );
  NAND2_X1 U94 ( .A1(n12), .A2(IN5[19]), .ZN(n102) );
  NAND4_X1 U95 ( .A1(n105), .A2(n104), .A3(n103), .A4(n102), .ZN(Y[19]) );
  AOI22_X1 U96 ( .A1(n10), .A2(IN0[1]), .B1(n9), .B2(IN1[1]), .ZN(n109) );
  AOI22_X1 U97 ( .A1(n8), .A2(IN2[1]), .B1(n7), .B2(IN3[1]), .ZN(n108) );
  AOI22_X1 U98 ( .A1(n6), .A2(IN6[1]), .B1(n11), .B2(IN4[1]), .ZN(n107) );
  NAND2_X1 U99 ( .A1(n12), .A2(IN5[1]), .ZN(n106) );
  NAND4_X1 U100 ( .A1(n109), .A2(n108), .A3(n107), .A4(n106), .ZN(Y[1]) );
  AOI22_X1 U101 ( .A1(n10), .A2(IN0[20]), .B1(n9), .B2(IN1[20]), .ZN(n113) );
  AOI22_X1 U102 ( .A1(n8), .A2(IN2[20]), .B1(n7), .B2(IN3[20]), .ZN(n112) );
  AOI22_X1 U103 ( .A1(n6), .A2(IN6[20]), .B1(n11), .B2(IN4[20]), .ZN(n111) );
  NAND2_X1 U104 ( .A1(n12), .A2(IN5[20]), .ZN(n110) );
  NAND4_X1 U105 ( .A1(n113), .A2(n112), .A3(n111), .A4(n110), .ZN(Y[20]) );
  AOI22_X1 U106 ( .A1(n10), .A2(IN0[21]), .B1(n9), .B2(IN1[21]), .ZN(n117) );
  AOI22_X1 U107 ( .A1(n8), .A2(IN2[21]), .B1(n7), .B2(IN3[21]), .ZN(n116) );
  AOI22_X1 U108 ( .A1(n6), .A2(IN6[21]), .B1(n11), .B2(IN4[21]), .ZN(n115) );
  NAND2_X1 U109 ( .A1(n12), .A2(IN5[21]), .ZN(n114) );
  NAND4_X1 U110 ( .A1(n117), .A2(n116), .A3(n115), .A4(n114), .ZN(Y[21]) );
  AOI22_X1 U111 ( .A1(n10), .A2(IN0[22]), .B1(n9), .B2(IN1[22]), .ZN(n121) );
  AOI22_X1 U112 ( .A1(n8), .A2(IN2[22]), .B1(n7), .B2(IN3[22]), .ZN(n120) );
  AOI22_X1 U113 ( .A1(n6), .A2(IN6[22]), .B1(n11), .B2(IN4[22]), .ZN(n119) );
  NAND2_X1 U114 ( .A1(n12), .A2(IN5[22]), .ZN(n118) );
  NAND4_X1 U115 ( .A1(n121), .A2(n120), .A3(n119), .A4(n118), .ZN(Y[22]) );
  AOI22_X1 U116 ( .A1(n10), .A2(IN0[23]), .B1(n9), .B2(IN1[23]), .ZN(n125) );
  AOI22_X1 U117 ( .A1(n8), .A2(IN2[23]), .B1(n7), .B2(IN3[23]), .ZN(n124) );
  AOI22_X1 U118 ( .A1(n6), .A2(IN6[23]), .B1(n11), .B2(IN4[23]), .ZN(n123) );
  NAND2_X1 U119 ( .A1(n12), .A2(IN5[23]), .ZN(n122) );
  NAND4_X1 U120 ( .A1(n125), .A2(n124), .A3(n123), .A4(n122), .ZN(Y[23]) );
  AOI22_X1 U121 ( .A1(n10), .A2(IN0[24]), .B1(n9), .B2(IN1[24]), .ZN(n129) );
  AOI22_X1 U122 ( .A1(n8), .A2(IN2[24]), .B1(n7), .B2(IN3[24]), .ZN(n128) );
  AOI22_X1 U123 ( .A1(n6), .A2(IN6[24]), .B1(n11), .B2(IN4[24]), .ZN(n127) );
  NAND2_X1 U124 ( .A1(n12), .A2(IN5[24]), .ZN(n126) );
  NAND4_X1 U125 ( .A1(n129), .A2(n128), .A3(n127), .A4(n126), .ZN(Y[24]) );
  AOI22_X1 U126 ( .A1(n10), .A2(IN0[25]), .B1(n9), .B2(IN1[25]), .ZN(n133) );
  AOI22_X1 U127 ( .A1(n8), .A2(IN2[25]), .B1(n7), .B2(IN3[25]), .ZN(n132) );
  AOI22_X1 U128 ( .A1(n6), .A2(IN6[25]), .B1(n11), .B2(IN4[25]), .ZN(n131) );
  NAND2_X1 U129 ( .A1(n12), .A2(IN5[25]), .ZN(n130) );
  NAND4_X1 U130 ( .A1(n133), .A2(n132), .A3(n131), .A4(n130), .ZN(Y[25]) );
  AOI22_X1 U131 ( .A1(n10), .A2(IN0[26]), .B1(n9), .B2(IN1[26]), .ZN(n137) );
  AOI22_X1 U132 ( .A1(n8), .A2(IN2[26]), .B1(n7), .B2(IN3[26]), .ZN(n136) );
  AOI22_X1 U133 ( .A1(n6), .A2(IN6[26]), .B1(n11), .B2(IN4[26]), .ZN(n135) );
  NAND2_X1 U134 ( .A1(n12), .A2(IN5[26]), .ZN(n134) );
  NAND4_X1 U135 ( .A1(n137), .A2(n136), .A3(n135), .A4(n134), .ZN(Y[26]) );
  AOI22_X1 U136 ( .A1(n10), .A2(IN0[27]), .B1(n9), .B2(IN1[27]), .ZN(n141) );
  AOI22_X1 U137 ( .A1(n8), .A2(IN2[27]), .B1(n7), .B2(IN3[27]), .ZN(n140) );
  AOI22_X1 U138 ( .A1(n6), .A2(IN6[27]), .B1(n11), .B2(IN4[27]), .ZN(n139) );
  NAND2_X1 U139 ( .A1(n12), .A2(IN5[27]), .ZN(n138) );
  NAND4_X1 U140 ( .A1(n141), .A2(n140), .A3(n139), .A4(n138), .ZN(Y[27]) );
  AOI22_X1 U141 ( .A1(n10), .A2(IN0[28]), .B1(n9), .B2(IN1[28]), .ZN(n145) );
  AOI22_X1 U142 ( .A1(n8), .A2(IN2[28]), .B1(n7), .B2(IN3[28]), .ZN(n144) );
  AOI22_X1 U143 ( .A1(n6), .A2(IN6[28]), .B1(n11), .B2(IN4[28]), .ZN(n143) );
  NAND2_X1 U144 ( .A1(n12), .A2(IN5[28]), .ZN(n142) );
  NAND4_X1 U145 ( .A1(n145), .A2(n144), .A3(n143), .A4(n142), .ZN(Y[28]) );
  AOI22_X1 U146 ( .A1(n10), .A2(IN0[29]), .B1(n9), .B2(IN1[29]), .ZN(n149) );
  AOI22_X1 U147 ( .A1(n8), .A2(IN2[29]), .B1(n7), .B2(IN3[29]), .ZN(n148) );
  AOI22_X1 U148 ( .A1(n6), .A2(IN6[29]), .B1(n11), .B2(IN4[29]), .ZN(n147) );
  NAND2_X1 U149 ( .A1(n12), .A2(IN5[29]), .ZN(n146) );
  NAND4_X1 U150 ( .A1(n149), .A2(n148), .A3(n147), .A4(n146), .ZN(Y[29]) );
  AOI22_X1 U151 ( .A1(n10), .A2(IN0[2]), .B1(n9), .B2(IN1[2]), .ZN(n153) );
  AOI22_X1 U152 ( .A1(n8), .A2(IN2[2]), .B1(n7), .B2(IN3[2]), .ZN(n152) );
  AOI22_X1 U153 ( .A1(n6), .A2(IN6[2]), .B1(n11), .B2(IN4[2]), .ZN(n151) );
  NAND2_X1 U154 ( .A1(n12), .A2(IN5[2]), .ZN(n150) );
  NAND4_X1 U155 ( .A1(n153), .A2(n152), .A3(n151), .A4(n150), .ZN(Y[2]) );
  AOI22_X1 U156 ( .A1(n8), .A2(IN2[31]), .B1(n7), .B2(IN3[31]), .ZN(n156) );
  AOI22_X1 U157 ( .A1(n6), .A2(IN6[31]), .B1(n11), .B2(IN4[31]), .ZN(n155) );
  NAND2_X1 U158 ( .A1(n12), .A2(IN5[31]), .ZN(n154) );
  AOI22_X1 U159 ( .A1(n10), .A2(IN0[3]), .B1(n9), .B2(IN1[3]), .ZN(n160) );
  AOI22_X1 U160 ( .A1(n8), .A2(IN2[3]), .B1(n7), .B2(IN3[3]), .ZN(n159) );
  AOI22_X1 U161 ( .A1(n6), .A2(IN6[3]), .B1(n11), .B2(IN4[3]), .ZN(n158) );
  NAND2_X1 U162 ( .A1(n12), .A2(IN5[3]), .ZN(n157) );
  NAND4_X1 U163 ( .A1(n160), .A2(n159), .A3(n158), .A4(n157), .ZN(Y[3]) );
  AOI22_X1 U164 ( .A1(n10), .A2(IN0[4]), .B1(n9), .B2(IN1[4]), .ZN(n164) );
  AOI22_X1 U165 ( .A1(n8), .A2(IN2[4]), .B1(n7), .B2(IN3[4]), .ZN(n163) );
  AOI22_X1 U166 ( .A1(n6), .A2(IN6[4]), .B1(n11), .B2(IN4[4]), .ZN(n162) );
  NAND2_X1 U167 ( .A1(n12), .A2(IN5[4]), .ZN(n161) );
  NAND4_X1 U168 ( .A1(n164), .A2(n163), .A3(n162), .A4(n161), .ZN(Y[4]) );
  AOI22_X1 U169 ( .A1(n10), .A2(IN0[5]), .B1(n9), .B2(IN1[5]), .ZN(n168) );
  AOI22_X1 U170 ( .A1(n8), .A2(IN2[5]), .B1(n7), .B2(IN3[5]), .ZN(n167) );
  AOI22_X1 U171 ( .A1(n6), .A2(IN6[5]), .B1(n11), .B2(IN4[5]), .ZN(n166) );
  NAND2_X1 U172 ( .A1(n12), .A2(IN5[5]), .ZN(n165) );
  NAND4_X1 U173 ( .A1(n168), .A2(n167), .A3(n166), .A4(n165), .ZN(Y[5]) );
  AOI22_X1 U174 ( .A1(n10), .A2(IN0[6]), .B1(n9), .B2(IN1[6]), .ZN(n172) );
  AOI22_X1 U175 ( .A1(n8), .A2(IN2[6]), .B1(n7), .B2(IN3[6]), .ZN(n171) );
  AOI22_X1 U176 ( .A1(n6), .A2(IN6[6]), .B1(n11), .B2(IN4[6]), .ZN(n170) );
  NAND2_X1 U177 ( .A1(n12), .A2(IN5[6]), .ZN(n169) );
  NAND4_X1 U178 ( .A1(n172), .A2(n171), .A3(n170), .A4(n169), .ZN(Y[6]) );
  AOI22_X1 U179 ( .A1(n8), .A2(IN2[7]), .B1(n7), .B2(IN3[7]), .ZN(n175) );
  AOI22_X1 U180 ( .A1(n6), .A2(IN6[7]), .B1(n11), .B2(IN4[7]), .ZN(n174) );
  NAND2_X1 U181 ( .A1(n12), .A2(IN5[7]), .ZN(n173) );
  AOI22_X1 U182 ( .A1(n10), .A2(IN0[8]), .B1(n9), .B2(IN1[8]), .ZN(n179) );
  AOI22_X1 U183 ( .A1(n8), .A2(IN2[8]), .B1(n7), .B2(IN3[8]), .ZN(n178) );
  AOI22_X1 U184 ( .A1(n6), .A2(IN6[8]), .B1(n11), .B2(IN4[8]), .ZN(n177) );
  NAND2_X1 U185 ( .A1(n12), .A2(IN5[8]), .ZN(n176) );
  NAND4_X1 U186 ( .A1(n179), .A2(n178), .A3(n177), .A4(n176), .ZN(Y[8]) );
  AOI22_X1 U187 ( .A1(n8), .A2(IN2[9]), .B1(n7), .B2(IN3[9]), .ZN(n189) );
  AOI22_X1 U188 ( .A1(n6), .A2(IN6[9]), .B1(n11), .B2(IN4[9]), .ZN(n188) );
  NAND2_X1 U189 ( .A1(n12), .A2(IN5[9]), .ZN(n187) );
endmodule


module MUX_8to1_N32_3 ( IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, SEL, Y );
  input [31:0] IN0;
  input [31:0] IN1;
  input [31:0] IN2;
  input [31:0] IN3;
  input [31:0] IN4;
  input [31:0] IN5;
  input [31:0] IN6;
  input [31:0] IN7;
  input [2:0] SEL;
  output [31:0] Y;
  wire   n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177;

  BUF_X2 U1 ( .A(n171), .Z(n35) );
  BUF_X2 U2 ( .A(n172), .Z(n34) );
  BUF_X2 U3 ( .A(n173), .Z(n33) );
  BUF_X2 U4 ( .A(n170), .Z(n36) );
  BUF_X2 U5 ( .A(n169), .Z(n37) );
  BUF_X2 U6 ( .A(n168), .Z(n38) );
  BUF_X2 U7 ( .A(n167), .Z(n39) );
  INV_X1 U8 ( .A(SEL[2]), .ZN(n41) );
  NOR3_X1 U9 ( .A1(SEL[2]), .A2(SEL[0]), .A3(SEL[1]), .ZN(n168) );
  INV_X1 U10 ( .A(SEL[0]), .ZN(n42) );
  NOR3_X1 U11 ( .A1(SEL[2]), .A2(SEL[1]), .A3(n42), .ZN(n167) );
  AOI22_X1 U12 ( .A1(n38), .A2(IN0[0]), .B1(n39), .B2(IN1[0]), .ZN(n46) );
  INV_X1 U13 ( .A(SEL[1]), .ZN(n40) );
  NOR3_X1 U14 ( .A1(SEL[2]), .A2(SEL[0]), .A3(n40), .ZN(n170) );
  NOR3_X1 U15 ( .A1(SEL[2]), .A2(n42), .A3(n40), .ZN(n169) );
  AOI22_X1 U16 ( .A1(n36), .A2(IN2[0]), .B1(n37), .B2(IN3[0]), .ZN(n45) );
  NOR3_X1 U17 ( .A1(SEL[0]), .A2(n41), .A3(n40), .ZN(n172) );
  NOR3_X1 U18 ( .A1(SEL[0]), .A2(SEL[1]), .A3(n41), .ZN(n171) );
  AOI22_X1 U19 ( .A1(n34), .A2(IN6[0]), .B1(n35), .B2(IN4[0]), .ZN(n44) );
  NOR3_X1 U20 ( .A1(SEL[1]), .A2(n42), .A3(n41), .ZN(n173) );
  NAND2_X1 U21 ( .A1(n33), .A2(IN5[0]), .ZN(n43) );
  NAND4_X1 U22 ( .A1(n46), .A2(n45), .A3(n44), .A4(n43), .ZN(Y[0]) );
  AOI22_X1 U23 ( .A1(n38), .A2(IN0[10]), .B1(n39), .B2(IN1[10]), .ZN(n50) );
  AOI22_X1 U24 ( .A1(n36), .A2(IN2[10]), .B1(n37), .B2(IN3[10]), .ZN(n49) );
  AOI22_X1 U25 ( .A1(n34), .A2(IN6[10]), .B1(n35), .B2(IN4[10]), .ZN(n48) );
  NAND2_X1 U26 ( .A1(n33), .A2(IN5[10]), .ZN(n47) );
  NAND4_X1 U27 ( .A1(n50), .A2(n49), .A3(n48), .A4(n47), .ZN(Y[10]) );
  AOI22_X1 U28 ( .A1(n38), .A2(IN0[11]), .B1(n39), .B2(IN1[11]), .ZN(n54) );
  AOI22_X1 U29 ( .A1(n36), .A2(IN2[11]), .B1(n37), .B2(IN3[11]), .ZN(n53) );
  AOI22_X1 U30 ( .A1(n34), .A2(IN6[11]), .B1(n35), .B2(IN4[11]), .ZN(n52) );
  NAND2_X1 U31 ( .A1(n33), .A2(IN5[11]), .ZN(n51) );
  NAND4_X1 U32 ( .A1(n54), .A2(n53), .A3(n52), .A4(n51), .ZN(Y[11]) );
  AOI22_X1 U33 ( .A1(n38), .A2(IN0[12]), .B1(n39), .B2(IN1[12]), .ZN(n58) );
  AOI22_X1 U34 ( .A1(n36), .A2(IN2[12]), .B1(n37), .B2(IN3[12]), .ZN(n57) );
  AOI22_X1 U35 ( .A1(n34), .A2(IN6[12]), .B1(n35), .B2(IN4[12]), .ZN(n56) );
  NAND2_X1 U36 ( .A1(n33), .A2(IN5[12]), .ZN(n55) );
  NAND4_X1 U37 ( .A1(n58), .A2(n57), .A3(n56), .A4(n55), .ZN(Y[12]) );
  AOI22_X1 U38 ( .A1(n38), .A2(IN0[13]), .B1(n39), .B2(IN1[13]), .ZN(n62) );
  AOI22_X1 U39 ( .A1(n36), .A2(IN2[13]), .B1(n37), .B2(IN3[13]), .ZN(n61) );
  AOI22_X1 U40 ( .A1(n34), .A2(IN6[13]), .B1(n35), .B2(IN4[13]), .ZN(n60) );
  NAND2_X1 U41 ( .A1(n33), .A2(IN5[13]), .ZN(n59) );
  NAND4_X1 U42 ( .A1(n62), .A2(n61), .A3(n60), .A4(n59), .ZN(Y[13]) );
  AOI22_X1 U43 ( .A1(n38), .A2(IN0[14]), .B1(n39), .B2(IN1[14]), .ZN(n66) );
  AOI22_X1 U44 ( .A1(n36), .A2(IN2[14]), .B1(n37), .B2(IN3[14]), .ZN(n65) );
  AOI22_X1 U45 ( .A1(n34), .A2(IN6[14]), .B1(n35), .B2(IN4[14]), .ZN(n64) );
  NAND2_X1 U46 ( .A1(n33), .A2(IN5[14]), .ZN(n63) );
  NAND4_X1 U47 ( .A1(n66), .A2(n65), .A3(n64), .A4(n63), .ZN(Y[14]) );
  AOI22_X1 U48 ( .A1(n38), .A2(IN0[15]), .B1(n39), .B2(IN1[15]), .ZN(n70) );
  AOI22_X1 U49 ( .A1(n36), .A2(IN2[15]), .B1(n37), .B2(IN3[15]), .ZN(n69) );
  AOI22_X1 U50 ( .A1(n34), .A2(IN6[15]), .B1(n35), .B2(IN4[15]), .ZN(n68) );
  NAND2_X1 U51 ( .A1(n33), .A2(IN5[15]), .ZN(n67) );
  NAND4_X1 U52 ( .A1(n70), .A2(n69), .A3(n68), .A4(n67), .ZN(Y[15]) );
  AOI22_X1 U53 ( .A1(n38), .A2(IN0[16]), .B1(n39), .B2(IN1[16]), .ZN(n74) );
  AOI22_X1 U54 ( .A1(n36), .A2(IN2[16]), .B1(n37), .B2(IN3[16]), .ZN(n73) );
  AOI22_X1 U55 ( .A1(n34), .A2(IN6[16]), .B1(n35), .B2(IN4[16]), .ZN(n72) );
  NAND2_X1 U56 ( .A1(n33), .A2(IN5[16]), .ZN(n71) );
  NAND4_X1 U57 ( .A1(n74), .A2(n73), .A3(n72), .A4(n71), .ZN(Y[16]) );
  AOI22_X1 U58 ( .A1(n38), .A2(IN0[17]), .B1(n39), .B2(IN1[17]), .ZN(n78) );
  AOI22_X1 U59 ( .A1(n36), .A2(IN2[17]), .B1(n37), .B2(IN3[17]), .ZN(n77) );
  AOI22_X1 U60 ( .A1(n34), .A2(IN6[17]), .B1(n35), .B2(IN4[17]), .ZN(n76) );
  NAND2_X1 U61 ( .A1(n33), .A2(IN5[17]), .ZN(n75) );
  NAND4_X1 U62 ( .A1(n78), .A2(n77), .A3(n76), .A4(n75), .ZN(Y[17]) );
  AOI22_X1 U63 ( .A1(n38), .A2(IN0[18]), .B1(n39), .B2(IN1[18]), .ZN(n82) );
  AOI22_X1 U64 ( .A1(n36), .A2(IN2[18]), .B1(n37), .B2(IN3[18]), .ZN(n81) );
  AOI22_X1 U65 ( .A1(n34), .A2(IN6[18]), .B1(n35), .B2(IN4[18]), .ZN(n80) );
  NAND2_X1 U66 ( .A1(n33), .A2(IN5[18]), .ZN(n79) );
  NAND4_X1 U67 ( .A1(n82), .A2(n81), .A3(n80), .A4(n79), .ZN(Y[18]) );
  AOI22_X1 U68 ( .A1(n38), .A2(IN0[19]), .B1(n39), .B2(IN1[19]), .ZN(n86) );
  AOI22_X1 U69 ( .A1(n36), .A2(IN2[19]), .B1(n37), .B2(IN3[19]), .ZN(n85) );
  AOI22_X1 U70 ( .A1(n34), .A2(IN6[19]), .B1(n35), .B2(IN4[19]), .ZN(n84) );
  NAND2_X1 U71 ( .A1(n33), .A2(IN5[19]), .ZN(n83) );
  NAND4_X1 U72 ( .A1(n86), .A2(n85), .A3(n84), .A4(n83), .ZN(Y[19]) );
  AOI22_X1 U73 ( .A1(n38), .A2(IN0[1]), .B1(n39), .B2(IN1[1]), .ZN(n90) );
  AOI22_X1 U74 ( .A1(n36), .A2(IN2[1]), .B1(n37), .B2(IN3[1]), .ZN(n89) );
  AOI22_X1 U75 ( .A1(n34), .A2(IN6[1]), .B1(n35), .B2(IN4[1]), .ZN(n88) );
  NAND2_X1 U76 ( .A1(n33), .A2(IN5[1]), .ZN(n87) );
  NAND4_X1 U77 ( .A1(n90), .A2(n89), .A3(n88), .A4(n87), .ZN(Y[1]) );
  AOI22_X1 U78 ( .A1(n38), .A2(IN0[20]), .B1(n39), .B2(IN1[20]), .ZN(n94) );
  AOI22_X1 U79 ( .A1(n36), .A2(IN2[20]), .B1(n37), .B2(IN3[20]), .ZN(n93) );
  AOI22_X1 U80 ( .A1(n34), .A2(IN6[20]), .B1(n35), .B2(IN4[20]), .ZN(n92) );
  NAND2_X1 U81 ( .A1(n33), .A2(IN5[20]), .ZN(n91) );
  NAND4_X1 U82 ( .A1(n94), .A2(n93), .A3(n92), .A4(n91), .ZN(Y[20]) );
  AOI22_X1 U83 ( .A1(n38), .A2(IN0[21]), .B1(n39), .B2(IN1[21]), .ZN(n98) );
  AOI22_X1 U84 ( .A1(n36), .A2(IN2[21]), .B1(n37), .B2(IN3[21]), .ZN(n97) );
  AOI22_X1 U85 ( .A1(n34), .A2(IN6[21]), .B1(n35), .B2(IN4[21]), .ZN(n96) );
  NAND2_X1 U86 ( .A1(n33), .A2(IN5[21]), .ZN(n95) );
  NAND4_X1 U87 ( .A1(n98), .A2(n97), .A3(n96), .A4(n95), .ZN(Y[21]) );
  AOI22_X1 U88 ( .A1(n38), .A2(IN0[22]), .B1(n39), .B2(IN1[22]), .ZN(n102) );
  AOI22_X1 U89 ( .A1(n36), .A2(IN2[22]), .B1(n37), .B2(IN3[22]), .ZN(n101) );
  AOI22_X1 U90 ( .A1(n34), .A2(IN6[22]), .B1(n35), .B2(IN4[22]), .ZN(n100) );
  NAND2_X1 U91 ( .A1(n33), .A2(IN5[22]), .ZN(n99) );
  NAND4_X1 U92 ( .A1(n102), .A2(n101), .A3(n100), .A4(n99), .ZN(Y[22]) );
  AOI22_X1 U93 ( .A1(n38), .A2(IN0[23]), .B1(n39), .B2(IN1[23]), .ZN(n106) );
  AOI22_X1 U94 ( .A1(n36), .A2(IN2[23]), .B1(n37), .B2(IN3[23]), .ZN(n105) );
  AOI22_X1 U95 ( .A1(n34), .A2(IN6[23]), .B1(n35), .B2(IN4[23]), .ZN(n104) );
  NAND2_X1 U96 ( .A1(n33), .A2(IN5[23]), .ZN(n103) );
  NAND4_X1 U97 ( .A1(n106), .A2(n105), .A3(n104), .A4(n103), .ZN(Y[23]) );
  AOI22_X1 U98 ( .A1(n38), .A2(IN0[24]), .B1(n39), .B2(IN1[24]), .ZN(n110) );
  AOI22_X1 U99 ( .A1(n36), .A2(IN2[24]), .B1(n37), .B2(IN3[24]), .ZN(n109) );
  AOI22_X1 U100 ( .A1(n34), .A2(IN6[24]), .B1(n35), .B2(IN4[24]), .ZN(n108) );
  NAND2_X1 U101 ( .A1(n33), .A2(IN5[24]), .ZN(n107) );
  NAND4_X1 U102 ( .A1(n110), .A2(n109), .A3(n108), .A4(n107), .ZN(Y[24]) );
  AOI22_X1 U103 ( .A1(n38), .A2(IN0[25]), .B1(n39), .B2(IN1[25]), .ZN(n114) );
  AOI22_X1 U104 ( .A1(n36), .A2(IN2[25]), .B1(n37), .B2(IN3[25]), .ZN(n113) );
  AOI22_X1 U105 ( .A1(n34), .A2(IN6[25]), .B1(n35), .B2(IN4[25]), .ZN(n112) );
  NAND2_X1 U106 ( .A1(n33), .A2(IN5[25]), .ZN(n111) );
  NAND4_X1 U107 ( .A1(n114), .A2(n113), .A3(n112), .A4(n111), .ZN(Y[25]) );
  AOI22_X1 U108 ( .A1(n38), .A2(IN0[26]), .B1(n39), .B2(IN1[26]), .ZN(n118) );
  AOI22_X1 U109 ( .A1(n36), .A2(IN2[26]), .B1(n37), .B2(IN3[26]), .ZN(n117) );
  AOI22_X1 U110 ( .A1(n34), .A2(IN6[26]), .B1(n35), .B2(IN4[26]), .ZN(n116) );
  NAND2_X1 U111 ( .A1(n33), .A2(IN5[26]), .ZN(n115) );
  NAND4_X1 U112 ( .A1(n118), .A2(n117), .A3(n116), .A4(n115), .ZN(Y[26]) );
  AOI22_X1 U113 ( .A1(n38), .A2(IN0[27]), .B1(n39), .B2(IN1[27]), .ZN(n122) );
  AOI22_X1 U114 ( .A1(n36), .A2(IN2[27]), .B1(n37), .B2(IN3[27]), .ZN(n121) );
  AOI22_X1 U115 ( .A1(n34), .A2(IN6[27]), .B1(n35), .B2(IN4[27]), .ZN(n120) );
  NAND2_X1 U116 ( .A1(n33), .A2(IN5[27]), .ZN(n119) );
  NAND4_X1 U117 ( .A1(n122), .A2(n121), .A3(n120), .A4(n119), .ZN(Y[27]) );
  AOI22_X1 U118 ( .A1(n38), .A2(IN0[28]), .B1(n39), .B2(IN1[28]), .ZN(n126) );
  AOI22_X1 U119 ( .A1(n36), .A2(IN2[28]), .B1(n37), .B2(IN3[28]), .ZN(n125) );
  AOI22_X1 U120 ( .A1(n34), .A2(IN6[28]), .B1(n35), .B2(IN4[28]), .ZN(n124) );
  NAND2_X1 U121 ( .A1(n33), .A2(IN5[28]), .ZN(n123) );
  NAND4_X1 U122 ( .A1(n126), .A2(n125), .A3(n124), .A4(n123), .ZN(Y[28]) );
  AOI22_X1 U123 ( .A1(n38), .A2(IN0[29]), .B1(n39), .B2(IN1[29]), .ZN(n130) );
  AOI22_X1 U124 ( .A1(n36), .A2(IN2[29]), .B1(n37), .B2(IN3[29]), .ZN(n129) );
  AOI22_X1 U125 ( .A1(n34), .A2(IN6[29]), .B1(n35), .B2(IN4[29]), .ZN(n128) );
  NAND2_X1 U126 ( .A1(n33), .A2(IN5[29]), .ZN(n127) );
  NAND4_X1 U127 ( .A1(n130), .A2(n129), .A3(n128), .A4(n127), .ZN(Y[29]) );
  AOI22_X1 U128 ( .A1(n38), .A2(IN0[2]), .B1(n39), .B2(IN1[2]), .ZN(n134) );
  AOI22_X1 U129 ( .A1(n36), .A2(IN2[2]), .B1(n37), .B2(IN3[2]), .ZN(n133) );
  AOI22_X1 U130 ( .A1(n34), .A2(IN6[2]), .B1(n35), .B2(IN4[2]), .ZN(n132) );
  NAND2_X1 U131 ( .A1(n33), .A2(IN5[2]), .ZN(n131) );
  NAND4_X1 U132 ( .A1(n134), .A2(n133), .A3(n132), .A4(n131), .ZN(Y[2]) );
  AOI22_X1 U133 ( .A1(n38), .A2(IN0[30]), .B1(n39), .B2(IN1[30]), .ZN(n138) );
  AOI22_X1 U134 ( .A1(n36), .A2(IN2[30]), .B1(n37), .B2(IN3[30]), .ZN(n137) );
  AOI22_X1 U135 ( .A1(n34), .A2(IN6[30]), .B1(n35), .B2(IN4[30]), .ZN(n136) );
  NAND2_X1 U136 ( .A1(n33), .A2(IN5[30]), .ZN(n135) );
  NAND4_X1 U137 ( .A1(n138), .A2(n137), .A3(n136), .A4(n135), .ZN(Y[30]) );
  AOI22_X1 U138 ( .A1(n38), .A2(IN0[31]), .B1(n39), .B2(IN1[31]), .ZN(n142) );
  AOI22_X1 U139 ( .A1(n36), .A2(IN2[31]), .B1(n37), .B2(IN3[31]), .ZN(n141) );
  AOI22_X1 U140 ( .A1(n34), .A2(IN6[31]), .B1(n35), .B2(IN4[31]), .ZN(n140) );
  NAND2_X1 U141 ( .A1(n33), .A2(IN5[31]), .ZN(n139) );
  NAND4_X1 U142 ( .A1(n142), .A2(n141), .A3(n140), .A4(n139), .ZN(Y[31]) );
  AOI22_X1 U143 ( .A1(n38), .A2(IN0[3]), .B1(n39), .B2(IN1[3]), .ZN(n146) );
  AOI22_X1 U144 ( .A1(n36), .A2(IN2[3]), .B1(n37), .B2(IN3[3]), .ZN(n145) );
  AOI22_X1 U145 ( .A1(n34), .A2(IN6[3]), .B1(n35), .B2(IN4[3]), .ZN(n144) );
  NAND2_X1 U146 ( .A1(n33), .A2(IN5[3]), .ZN(n143) );
  NAND4_X1 U147 ( .A1(n146), .A2(n145), .A3(n144), .A4(n143), .ZN(Y[3]) );
  AOI22_X1 U148 ( .A1(n38), .A2(IN0[4]), .B1(n39), .B2(IN1[4]), .ZN(n150) );
  AOI22_X1 U149 ( .A1(n36), .A2(IN2[4]), .B1(n37), .B2(IN3[4]), .ZN(n149) );
  AOI22_X1 U150 ( .A1(n34), .A2(IN6[4]), .B1(n35), .B2(IN4[4]), .ZN(n148) );
  NAND2_X1 U151 ( .A1(n33), .A2(IN5[4]), .ZN(n147) );
  NAND4_X1 U152 ( .A1(n150), .A2(n149), .A3(n148), .A4(n147), .ZN(Y[4]) );
  AOI22_X1 U153 ( .A1(n168), .A2(IN0[5]), .B1(n39), .B2(IN1[5]), .ZN(n154) );
  AOI22_X1 U154 ( .A1(n36), .A2(IN2[5]), .B1(n37), .B2(IN3[5]), .ZN(n153) );
  AOI22_X1 U155 ( .A1(n34), .A2(IN6[5]), .B1(n35), .B2(IN4[5]), .ZN(n152) );
  NAND2_X1 U156 ( .A1(n33), .A2(IN5[5]), .ZN(n151) );
  NAND4_X1 U157 ( .A1(n154), .A2(n153), .A3(n152), .A4(n151), .ZN(Y[5]) );
  AOI22_X1 U158 ( .A1(n38), .A2(IN0[6]), .B1(n39), .B2(IN1[6]), .ZN(n158) );
  AOI22_X1 U159 ( .A1(n36), .A2(IN2[6]), .B1(n37), .B2(IN3[6]), .ZN(n157) );
  AOI22_X1 U160 ( .A1(n34), .A2(IN6[6]), .B1(n35), .B2(IN4[6]), .ZN(n156) );
  NAND2_X1 U161 ( .A1(n33), .A2(IN5[6]), .ZN(n155) );
  NAND4_X1 U162 ( .A1(n158), .A2(n157), .A3(n156), .A4(n155), .ZN(Y[6]) );
  AOI22_X1 U163 ( .A1(n38), .A2(IN0[7]), .B1(n39), .B2(IN1[7]), .ZN(n162) );
  AOI22_X1 U164 ( .A1(n36), .A2(IN2[7]), .B1(n37), .B2(IN3[7]), .ZN(n161) );
  AOI22_X1 U165 ( .A1(n34), .A2(IN6[7]), .B1(n35), .B2(IN4[7]), .ZN(n160) );
  NAND2_X1 U166 ( .A1(n33), .A2(IN5[7]), .ZN(n159) );
  NAND4_X1 U167 ( .A1(n162), .A2(n161), .A3(n160), .A4(n159), .ZN(Y[7]) );
  AOI22_X1 U168 ( .A1(n38), .A2(IN0[8]), .B1(n39), .B2(IN1[8]), .ZN(n166) );
  AOI22_X1 U169 ( .A1(n36), .A2(IN2[8]), .B1(n37), .B2(IN3[8]), .ZN(n165) );
  AOI22_X1 U170 ( .A1(n34), .A2(IN6[8]), .B1(n35), .B2(IN4[8]), .ZN(n164) );
  NAND2_X1 U171 ( .A1(n33), .A2(IN5[8]), .ZN(n163) );
  NAND4_X1 U172 ( .A1(n166), .A2(n165), .A3(n164), .A4(n163), .ZN(Y[8]) );
  AOI22_X1 U173 ( .A1(n38), .A2(IN0[9]), .B1(n39), .B2(IN1[9]), .ZN(n177) );
  AOI22_X1 U174 ( .A1(n36), .A2(IN2[9]), .B1(n37), .B2(IN3[9]), .ZN(n176) );
  AOI22_X1 U175 ( .A1(n34), .A2(IN6[9]), .B1(n35), .B2(IN4[9]), .ZN(n175) );
  NAND2_X1 U176 ( .A1(n33), .A2(IN5[9]), .ZN(n174) );
  NAND4_X1 U177 ( .A1(n177), .A2(n176), .A3(n175), .A4(n174), .ZN(Y[9]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_reg_N32_10 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18782, net18784, net18786, net18787, net18790, net18793;
  assign net18782 = EN;
  assign net18784 = CLK;
  assign ENCLK = net18786;
  assign net18793 = TE;

  DLL_X1 latch ( .D(net18787), .GN(net18784), .Q(net18790) );
  AND2_X1 main_gate ( .A1(net18790), .A2(net18784), .ZN(net18786) );
  OR2_X1 test_or ( .A1(net18782), .A2(net18793), .ZN(net18787) );
endmodule


module reg_N32_10 ( D, Q, EN, CLK, RST );
  input [31:0] D;
  output [31:0] Q;
  input EN, CLK, RST;
  wire   net18798;

  SNPS_CLOCK_GATE_HIGH_reg_N32_10 clk_gate_Q_reg ( .CLK(CLK), .EN(EN), .ENCLK(
        net18798), .TE(1'b0) );
  DFFR_X1 \Q_reg[31]  ( .D(D[31]), .CK(net18798), .RN(RST), .Q(Q[31]) );
  DFFR_X1 \Q_reg[30]  ( .D(D[30]), .CK(net18798), .RN(RST), .Q(Q[30]) );
  DFFR_X1 \Q_reg[29]  ( .D(D[29]), .CK(net18798), .RN(RST), .Q(Q[29]) );
  DFFR_X1 \Q_reg[28]  ( .D(D[28]), .CK(net18798), .RN(RST), .Q(Q[28]) );
  DFFR_X1 \Q_reg[27]  ( .D(D[27]), .CK(net18798), .RN(RST), .Q(Q[27]) );
  DFFR_X1 \Q_reg[26]  ( .D(D[26]), .CK(net18798), .RN(RST), .Q(Q[26]) );
  DFFR_X1 \Q_reg[25]  ( .D(D[25]), .CK(net18798), .RN(RST), .Q(Q[25]) );
  DFFR_X1 \Q_reg[24]  ( .D(D[24]), .CK(net18798), .RN(RST), .Q(Q[24]) );
  DFFR_X1 \Q_reg[23]  ( .D(D[23]), .CK(net18798), .RN(RST), .Q(Q[23]) );
  DFFR_X1 \Q_reg[22]  ( .D(D[22]), .CK(net18798), .RN(RST), .Q(Q[22]) );
  DFFR_X1 \Q_reg[21]  ( .D(D[21]), .CK(net18798), .RN(RST), .Q(Q[21]) );
  DFFR_X1 \Q_reg[20]  ( .D(D[20]), .CK(net18798), .RN(RST), .Q(Q[20]) );
  DFFR_X1 \Q_reg[19]  ( .D(D[19]), .CK(net18798), .RN(RST), .Q(Q[19]) );
  DFFR_X1 \Q_reg[18]  ( .D(D[18]), .CK(net18798), .RN(RST), .Q(Q[18]) );
  DFFR_X1 \Q_reg[17]  ( .D(D[17]), .CK(net18798), .RN(RST), .Q(Q[17]) );
  DFFR_X1 \Q_reg[16]  ( .D(D[16]), .CK(net18798), .RN(RST), .Q(Q[16]) );
  DFFR_X1 \Q_reg[15]  ( .D(D[15]), .CK(net18798), .RN(RST), .Q(Q[15]) );
  DFFR_X1 \Q_reg[14]  ( .D(D[14]), .CK(net18798), .RN(RST), .Q(Q[14]) );
  DFFR_X1 \Q_reg[13]  ( .D(D[13]), .CK(net18798), .RN(RST), .Q(Q[13]) );
  DFFR_X1 \Q_reg[12]  ( .D(D[12]), .CK(net18798), .RN(RST), .Q(Q[12]) );
  DFFR_X1 \Q_reg[11]  ( .D(D[11]), .CK(net18798), .RN(RST), .Q(Q[11]) );
  DFFR_X1 \Q_reg[10]  ( .D(D[10]), .CK(net18798), .RN(RST), .Q(Q[10]) );
  DFFR_X1 \Q_reg[9]  ( .D(D[9]), .CK(net18798), .RN(RST), .Q(Q[9]) );
  DFFR_X1 \Q_reg[8]  ( .D(D[8]), .CK(net18798), .RN(RST), .Q(Q[8]) );
  DFFR_X1 \Q_reg[7]  ( .D(D[7]), .CK(net18798), .RN(RST), .Q(Q[7]) );
  DFFR_X1 \Q_reg[6]  ( .D(D[6]), .CK(net18798), .RN(RST), .Q(Q[6]) );
  DFFR_X1 \Q_reg[5]  ( .D(D[5]), .CK(net18798), .RN(RST), .Q(Q[5]) );
  DFFR_X1 \Q_reg[4]  ( .D(D[4]), .CK(net18798), .RN(RST), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(D[3]), .CK(net18798), .RN(RST), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(D[2]), .CK(net18798), .RN(RST), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(D[1]), .CK(net18798), .RN(RST), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(D[0]), .CK(net18798), .RN(RST), .Q(Q[0]) );
endmodule


module MUX_4to1_N5 ( IN0, IN1, IN2, IN3, SEL, Y );
  input [4:0] IN0;
  input [4:0] IN1;
  input [4:0] IN2;
  input [4:0] IN3;
  input [1:0] SEL;
  output [4:0] Y;
  wire   n1, n2, n3, n4, n5, n6, n7, n8;

  INV_X1 U1 ( .A(SEL[0]), .ZN(n5) );
  NOR2_X1 U2 ( .A1(SEL[1]), .A2(n5), .ZN(n6) );
  AOI22_X1 U3 ( .A1(IN1[0]), .A2(n6), .B1(IN0[0]), .B2(n5), .ZN(n1) );
  NAND2_X1 U4 ( .A1(SEL[1]), .A2(n5), .ZN(n7) );
  NAND2_X1 U5 ( .A1(n1), .A2(n7), .ZN(Y[0]) );
  AOI22_X1 U6 ( .A1(IN1[1]), .A2(n6), .B1(IN0[1]), .B2(n5), .ZN(n2) );
  NAND2_X1 U7 ( .A1(n2), .A2(n7), .ZN(Y[1]) );
  AOI22_X1 U8 ( .A1(IN1[2]), .A2(n6), .B1(IN0[2]), .B2(n5), .ZN(n3) );
  NAND2_X1 U9 ( .A1(n3), .A2(n7), .ZN(Y[2]) );
  AOI22_X1 U10 ( .A1(IN1[3]), .A2(n6), .B1(IN0[3]), .B2(n5), .ZN(n4) );
  NAND2_X1 U11 ( .A1(n4), .A2(n7), .ZN(Y[3]) );
  AOI22_X1 U12 ( .A1(IN1[4]), .A2(n6), .B1(IN0[4]), .B2(n5), .ZN(n8) );
  NAND2_X1 U13 ( .A1(n8), .A2(n7), .ZN(Y[4]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_reg_N5_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18764, net18766, net18768, net18769, net18772, net18775;
  assign net18764 = EN;
  assign net18766 = CLK;
  assign ENCLK = net18768;
  assign net18775 = TE;

  DLL_X1 latch ( .D(net18769), .GN(net18766), .Q(net18772) );
  AND2_X1 main_gate ( .A1(net18772), .A2(net18766), .ZN(net18768) );
  OR2_X1 test_or ( .A1(net18764), .A2(net18775), .ZN(net18769) );
endmodule


module reg_N5_0 ( D, Q, EN, CLK, RST );
  input [4:0] D;
  output [4:0] Q;
  input EN, CLK, RST;
  wire   net18780;

  SNPS_CLOCK_GATE_HIGH_reg_N5_0 clk_gate_Q_reg ( .CLK(CLK), .EN(EN), .ENCLK(
        net18780), .TE(1'b0) );
  DFFR_X1 \Q_reg[4]  ( .D(D[4]), .CK(net18780), .RN(RST), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(D[3]), .CK(net18780), .RN(RST), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(D[2]), .CK(net18780), .RN(RST), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(D[1]), .CK(net18780), .RN(RST), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(D[0]), .CK(net18780), .RN(RST), .Q(Q[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_0 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18843, net18845, net18847, net18848, net18851, net18854;
  assign net18843 = EN;
  assign net18845 = CLK;
  assign ENCLK = net18847;
  assign net18854 = TE;

  DLL_X1 latch ( .D(net18848), .GN(net18845), .Q(net18851) );
  AND2_X1 main_gate ( .A1(net18851), .A2(net18845), .ZN(net18847) );
  OR2_X1 test_or ( .A1(net18843), .A2(net18854), .ZN(net18848) );
endmodule


module SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_30 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18843, net18845, net18847, net18848, net18851, net18854;
  assign net18843 = EN;
  assign net18845 = CLK;
  assign ENCLK = net18847;
  assign net18854 = TE;

  DLL_X1 latch ( .D(net18848), .GN(net18845), .Q(net18851) );
  AND2_X1 main_gate ( .A1(net18851), .A2(net18845), .ZN(net18847) );
  OR2_X1 test_or ( .A1(net18843), .A2(net18854), .ZN(net18848) );
endmodule


module SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_29 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18843, net18845, net18847, net18848, net18851, net18854;
  assign net18843 = EN;
  assign net18845 = CLK;
  assign ENCLK = net18847;
  assign net18854 = TE;

  DLL_X1 latch ( .D(net18848), .GN(net18845), .Q(net18851) );
  AND2_X1 main_gate ( .A1(net18851), .A2(net18845), .ZN(net18847) );
  OR2_X1 test_or ( .A1(net18843), .A2(net18854), .ZN(net18848) );
endmodule


module SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_28 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18843, net18845, net18847, net18848, net18851, net18854;
  assign net18843 = EN;
  assign net18845 = CLK;
  assign ENCLK = net18847;
  assign net18854 = TE;

  DLL_X1 latch ( .D(net18848), .GN(net18845), .Q(net18851) );
  AND2_X1 main_gate ( .A1(net18851), .A2(net18845), .ZN(net18847) );
  OR2_X1 test_or ( .A1(net18843), .A2(net18854), .ZN(net18848) );
endmodule


module SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_27 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18843, net18845, net18847, net18848, net18851, net18854;
  assign net18843 = EN;
  assign net18845 = CLK;
  assign ENCLK = net18847;
  assign net18854 = TE;

  DLL_X1 latch ( .D(net18848), .GN(net18845), .Q(net18851) );
  AND2_X1 main_gate ( .A1(net18851), .A2(net18845), .ZN(net18847) );
  OR2_X1 test_or ( .A1(net18843), .A2(net18854), .ZN(net18848) );
endmodule


module SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_26 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18843, net18845, net18847, net18848, net18851, net18854;
  assign net18843 = EN;
  assign net18845 = CLK;
  assign ENCLK = net18847;
  assign net18854 = TE;

  DLL_X1 latch ( .D(net18848), .GN(net18845), .Q(net18851) );
  AND2_X1 main_gate ( .A1(net18851), .A2(net18845), .ZN(net18847) );
  OR2_X1 test_or ( .A1(net18843), .A2(net18854), .ZN(net18848) );
endmodule


module SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_25 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18843, net18845, net18847, net18848, net18851, net18854;
  assign net18843 = EN;
  assign net18845 = CLK;
  assign ENCLK = net18847;
  assign net18854 = TE;

  DLL_X1 latch ( .D(net18848), .GN(net18845), .Q(net18851) );
  AND2_X1 main_gate ( .A1(net18851), .A2(net18845), .ZN(net18847) );
  OR2_X1 test_or ( .A1(net18843), .A2(net18854), .ZN(net18848) );
endmodule


module SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_24 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18843, net18845, net18847, net18848, net18851, net18854;
  assign net18843 = EN;
  assign net18845 = CLK;
  assign ENCLK = net18847;
  assign net18854 = TE;

  DLL_X1 latch ( .D(net18848), .GN(net18845), .Q(net18851) );
  AND2_X1 main_gate ( .A1(net18851), .A2(net18845), .ZN(net18847) );
  OR2_X1 test_or ( .A1(net18843), .A2(net18854), .ZN(net18848) );
endmodule


module SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_23 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18843, net18845, net18847, net18848, net18851, net18854;
  assign net18843 = EN;
  assign net18845 = CLK;
  assign ENCLK = net18847;
  assign net18854 = TE;

  DLL_X1 latch ( .D(net18848), .GN(net18845), .Q(net18851) );
  AND2_X1 main_gate ( .A1(net18851), .A2(net18845), .ZN(net18847) );
  OR2_X1 test_or ( .A1(net18843), .A2(net18854), .ZN(net18848) );
endmodule


module SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_22 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18843, net18845, net18847, net18848, net18851, net18854;
  assign net18843 = EN;
  assign net18845 = CLK;
  assign ENCLK = net18847;
  assign net18854 = TE;

  DLL_X1 latch ( .D(net18848), .GN(net18845), .Q(net18851) );
  AND2_X1 main_gate ( .A1(net18851), .A2(net18845), .ZN(net18847) );
  OR2_X1 test_or ( .A1(net18843), .A2(net18854), .ZN(net18848) );
endmodule


module SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_21 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18843, net18845, net18847, net18848, net18851, net18854;
  assign net18843 = EN;
  assign net18845 = CLK;
  assign ENCLK = net18847;
  assign net18854 = TE;

  DLL_X1 latch ( .D(net18848), .GN(net18845), .Q(net18851) );
  AND2_X1 main_gate ( .A1(net18851), .A2(net18845), .ZN(net18847) );
  OR2_X1 test_or ( .A1(net18843), .A2(net18854), .ZN(net18848) );
endmodule


module SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_20 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18843, net18845, net18847, net18848, net18851, net18854;
  assign net18843 = EN;
  assign net18845 = CLK;
  assign ENCLK = net18847;
  assign net18854 = TE;

  DLL_X1 latch ( .D(net18848), .GN(net18845), .Q(net18851) );
  AND2_X1 main_gate ( .A1(net18851), .A2(net18845), .ZN(net18847) );
  OR2_X1 test_or ( .A1(net18843), .A2(net18854), .ZN(net18848) );
endmodule


module SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_19 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18843, net18845, net18847, net18848, net18851, net18854;
  assign net18843 = EN;
  assign net18845 = CLK;
  assign ENCLK = net18847;
  assign net18854 = TE;

  DLL_X1 latch ( .D(net18848), .GN(net18845), .Q(net18851) );
  AND2_X1 main_gate ( .A1(net18851), .A2(net18845), .ZN(net18847) );
  OR2_X1 test_or ( .A1(net18843), .A2(net18854), .ZN(net18848) );
endmodule


module SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_18 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18843, net18845, net18847, net18848, net18851, net18854;
  assign net18843 = EN;
  assign net18845 = CLK;
  assign ENCLK = net18847;
  assign net18854 = TE;

  DLL_X1 latch ( .D(net18848), .GN(net18845), .Q(net18851) );
  AND2_X1 main_gate ( .A1(net18851), .A2(net18845), .ZN(net18847) );
  OR2_X1 test_or ( .A1(net18843), .A2(net18854), .ZN(net18848) );
endmodule


module SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_17 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18843, net18845, net18847, net18848, net18851, net18854;
  assign net18843 = EN;
  assign net18845 = CLK;
  assign ENCLK = net18847;
  assign net18854 = TE;

  DLL_X1 latch ( .D(net18848), .GN(net18845), .Q(net18851) );
  AND2_X1 main_gate ( .A1(net18851), .A2(net18845), .ZN(net18847) );
  OR2_X1 test_or ( .A1(net18843), .A2(net18854), .ZN(net18848) );
endmodule


module SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_16 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18843, net18845, net18847, net18848, net18851, net18854;
  assign net18843 = EN;
  assign net18845 = CLK;
  assign ENCLK = net18847;
  assign net18854 = TE;

  DLL_X1 latch ( .D(net18848), .GN(net18845), .Q(net18851) );
  AND2_X1 main_gate ( .A1(net18851), .A2(net18845), .ZN(net18847) );
  OR2_X1 test_or ( .A1(net18843), .A2(net18854), .ZN(net18848) );
endmodule


module SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_15 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18843, net18845, net18847, net18848, net18851, net18854;
  assign net18843 = EN;
  assign net18845 = CLK;
  assign ENCLK = net18847;
  assign net18854 = TE;

  DLL_X1 latch ( .D(net18848), .GN(net18845), .Q(net18851) );
  AND2_X1 main_gate ( .A1(net18851), .A2(net18845), .ZN(net18847) );
  OR2_X1 test_or ( .A1(net18843), .A2(net18854), .ZN(net18848) );
endmodule


module SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_14 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18843, net18845, net18847, net18848, net18851, net18854;
  assign net18843 = EN;
  assign net18845 = CLK;
  assign ENCLK = net18847;
  assign net18854 = TE;

  DLL_X1 latch ( .D(net18848), .GN(net18845), .Q(net18851) );
  AND2_X1 main_gate ( .A1(net18851), .A2(net18845), .ZN(net18847) );
  OR2_X1 test_or ( .A1(net18843), .A2(net18854), .ZN(net18848) );
endmodule


module SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_13 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18843, net18845, net18847, net18848, net18851, net18854;
  assign net18843 = EN;
  assign net18845 = CLK;
  assign ENCLK = net18847;
  assign net18854 = TE;

  DLL_X1 latch ( .D(net18848), .GN(net18845), .Q(net18851) );
  AND2_X1 main_gate ( .A1(net18851), .A2(net18845), .ZN(net18847) );
  OR2_X1 test_or ( .A1(net18843), .A2(net18854), .ZN(net18848) );
endmodule


module SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_12 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18843, net18845, net18847, net18848, net18851, net18854;
  assign net18843 = EN;
  assign net18845 = CLK;
  assign ENCLK = net18847;
  assign net18854 = TE;

  DLL_X1 latch ( .D(net18848), .GN(net18845), .Q(net18851) );
  AND2_X1 main_gate ( .A1(net18851), .A2(net18845), .ZN(net18847) );
  OR2_X1 test_or ( .A1(net18843), .A2(net18854), .ZN(net18848) );
endmodule


module SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_11 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18843, net18845, net18847, net18848, net18851, net18854;
  assign net18843 = EN;
  assign net18845 = CLK;
  assign ENCLK = net18847;
  assign net18854 = TE;

  DLL_X1 latch ( .D(net18848), .GN(net18845), .Q(net18851) );
  AND2_X1 main_gate ( .A1(net18851), .A2(net18845), .ZN(net18847) );
  OR2_X1 test_or ( .A1(net18843), .A2(net18854), .ZN(net18848) );
endmodule


module SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_10 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18843, net18845, net18847, net18848, net18851, net18854;
  assign net18843 = EN;
  assign net18845 = CLK;
  assign ENCLK = net18847;
  assign net18854 = TE;

  DLL_X1 latch ( .D(net18848), .GN(net18845), .Q(net18851) );
  AND2_X1 main_gate ( .A1(net18851), .A2(net18845), .ZN(net18847) );
  OR2_X1 test_or ( .A1(net18843), .A2(net18854), .ZN(net18848) );
endmodule


module SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_9 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18843, net18845, net18847, net18848, net18851, net18854;
  assign net18843 = EN;
  assign net18845 = CLK;
  assign ENCLK = net18847;
  assign net18854 = TE;

  DLL_X1 latch ( .D(net18848), .GN(net18845), .Q(net18851) );
  AND2_X1 main_gate ( .A1(net18851), .A2(net18845), .ZN(net18847) );
  OR2_X1 test_or ( .A1(net18843), .A2(net18854), .ZN(net18848) );
endmodule


module SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_8 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18843, net18845, net18847, net18848, net18851, net18854;
  assign net18843 = EN;
  assign net18845 = CLK;
  assign ENCLK = net18847;
  assign net18854 = TE;

  DLL_X1 latch ( .D(net18848), .GN(net18845), .Q(net18851) );
  AND2_X1 main_gate ( .A1(net18851), .A2(net18845), .ZN(net18847) );
  OR2_X1 test_or ( .A1(net18843), .A2(net18854), .ZN(net18848) );
endmodule


module SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_7 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18843, net18845, net18847, net18848, net18851, net18854;
  assign net18843 = EN;
  assign net18845 = CLK;
  assign ENCLK = net18847;
  assign net18854 = TE;

  DLL_X1 latch ( .D(net18848), .GN(net18845), .Q(net18851) );
  AND2_X1 main_gate ( .A1(net18851), .A2(net18845), .ZN(net18847) );
  OR2_X1 test_or ( .A1(net18843), .A2(net18854), .ZN(net18848) );
endmodule


module SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18843, net18845, net18847, net18848, net18851, net18854;
  assign net18843 = EN;
  assign net18845 = CLK;
  assign ENCLK = net18847;
  assign net18854 = TE;

  DLL_X1 latch ( .D(net18848), .GN(net18845), .Q(net18851) );
  AND2_X1 main_gate ( .A1(net18851), .A2(net18845), .ZN(net18847) );
  OR2_X1 test_or ( .A1(net18843), .A2(net18854), .ZN(net18848) );
endmodule


module SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18843, net18845, net18847, net18848, net18851, net18854;
  assign net18843 = EN;
  assign net18845 = CLK;
  assign ENCLK = net18847;
  assign net18854 = TE;

  DLL_X1 latch ( .D(net18848), .GN(net18845), .Q(net18851) );
  AND2_X1 main_gate ( .A1(net18851), .A2(net18845), .ZN(net18847) );
  OR2_X1 test_or ( .A1(net18843), .A2(net18854), .ZN(net18848) );
endmodule


module SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18843, net18845, net18847, net18848, net18851, net18854;
  assign net18843 = EN;
  assign net18845 = CLK;
  assign ENCLK = net18847;
  assign net18854 = TE;

  DLL_X1 latch ( .D(net18848), .GN(net18845), .Q(net18851) );
  AND2_X1 main_gate ( .A1(net18851), .A2(net18845), .ZN(net18847) );
  OR2_X1 test_or ( .A1(net18843), .A2(net18854), .ZN(net18848) );
endmodule


module SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18843, net18845, net18847, net18848, net18851, net18854;
  assign net18843 = EN;
  assign net18845 = CLK;
  assign ENCLK = net18847;
  assign net18854 = TE;

  DLL_X1 latch ( .D(net18848), .GN(net18845), .Q(net18851) );
  AND2_X1 main_gate ( .A1(net18851), .A2(net18845), .ZN(net18847) );
  OR2_X1 test_or ( .A1(net18843), .A2(net18854), .ZN(net18848) );
endmodule


module SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18843, net18845, net18847, net18848, net18851, net18854;
  assign net18843 = EN;
  assign net18845 = CLK;
  assign ENCLK = net18847;
  assign net18854 = TE;

  DLL_X1 latch ( .D(net18848), .GN(net18845), .Q(net18851) );
  AND2_X1 main_gate ( .A1(net18851), .A2(net18845), .ZN(net18847) );
  OR2_X1 test_or ( .A1(net18843), .A2(net18854), .ZN(net18848) );
endmodule


module SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18843, net18845, net18847, net18848, net18851, net18854;
  assign net18843 = EN;
  assign net18845 = CLK;
  assign ENCLK = net18847;
  assign net18854 = TE;

  DLL_X1 latch ( .D(net18848), .GN(net18845), .Q(net18851) );
  AND2_X1 main_gate ( .A1(net18851), .A2(net18845), .ZN(net18847) );
  OR2_X1 test_or ( .A1(net18843), .A2(net18854), .ZN(net18848) );
endmodule


module RF_N_bit32_N_reg32 ( CLK, RST, WR_EN, ADD_WR, ADD_RD1, ADD_RD2, DATA_IN, 
        OUT1, OUT2 );
  input [4:0] ADD_WR;
  input [4:0] ADD_RD1;
  input [4:0] ADD_RD2;
  input [31:0] DATA_IN;
  output [31:0] OUT1;
  output [31:0] OUT2;
  input CLK, RST, WR_EN;
  wire   \REGISTERS[1][31] , \REGISTERS[1][30] , \REGISTERS[1][29] ,
         \REGISTERS[1][28] , \REGISTERS[1][27] , \REGISTERS[1][26] ,
         \REGISTERS[1][25] , \REGISTERS[1][24] , \REGISTERS[1][23] ,
         \REGISTERS[1][22] , \REGISTERS[1][21] , \REGISTERS[1][20] ,
         \REGISTERS[1][19] , \REGISTERS[1][18] , \REGISTERS[1][17] ,
         \REGISTERS[1][16] , \REGISTERS[1][15] , \REGISTERS[1][14] ,
         \REGISTERS[1][13] , \REGISTERS[1][12] , \REGISTERS[1][11] ,
         \REGISTERS[1][10] , \REGISTERS[1][9] , \REGISTERS[1][8] ,
         \REGISTERS[1][7] , \REGISTERS[1][6] , \REGISTERS[1][5] ,
         \REGISTERS[1][4] , \REGISTERS[1][3] , \REGISTERS[1][2] ,
         \REGISTERS[1][1] , \REGISTERS[1][0] , \REGISTERS[2][31] ,
         \REGISTERS[2][30] , \REGISTERS[2][29] , \REGISTERS[2][28] ,
         \REGISTERS[2][27] , \REGISTERS[2][26] , \REGISTERS[2][25] ,
         \REGISTERS[2][24] , \REGISTERS[2][23] , \REGISTERS[2][22] ,
         \REGISTERS[2][21] , \REGISTERS[2][20] , \REGISTERS[2][19] ,
         \REGISTERS[2][18] , \REGISTERS[2][17] , \REGISTERS[2][16] ,
         \REGISTERS[2][15] , \REGISTERS[2][14] , \REGISTERS[2][13] ,
         \REGISTERS[2][12] , \REGISTERS[2][11] , \REGISTERS[2][10] ,
         \REGISTERS[2][9] , \REGISTERS[2][8] , \REGISTERS[2][7] ,
         \REGISTERS[2][6] , \REGISTERS[2][5] , \REGISTERS[2][4] ,
         \REGISTERS[2][3] , \REGISTERS[2][2] , \REGISTERS[2][1] ,
         \REGISTERS[2][0] , \REGISTERS[3][31] , \REGISTERS[3][30] ,
         \REGISTERS[3][29] , \REGISTERS[3][28] , \REGISTERS[3][27] ,
         \REGISTERS[3][26] , \REGISTERS[3][25] , \REGISTERS[3][24] ,
         \REGISTERS[3][23] , \REGISTERS[3][22] , \REGISTERS[3][21] ,
         \REGISTERS[3][20] , \REGISTERS[3][19] , \REGISTERS[3][18] ,
         \REGISTERS[3][17] , \REGISTERS[3][16] , \REGISTERS[3][15] ,
         \REGISTERS[3][14] , \REGISTERS[3][13] , \REGISTERS[3][12] ,
         \REGISTERS[3][11] , \REGISTERS[3][10] , \REGISTERS[3][9] ,
         \REGISTERS[3][8] , \REGISTERS[3][7] , \REGISTERS[3][6] ,
         \REGISTERS[3][5] , \REGISTERS[3][4] , \REGISTERS[3][3] ,
         \REGISTERS[3][2] , \REGISTERS[3][1] , \REGISTERS[3][0] ,
         \REGISTERS[4][31] , \REGISTERS[4][30] , \REGISTERS[4][29] ,
         \REGISTERS[4][28] , \REGISTERS[4][27] , \REGISTERS[4][26] ,
         \REGISTERS[4][25] , \REGISTERS[4][24] , \REGISTERS[4][23] ,
         \REGISTERS[4][22] , \REGISTERS[4][21] , \REGISTERS[4][20] ,
         \REGISTERS[4][19] , \REGISTERS[4][18] , \REGISTERS[4][17] ,
         \REGISTERS[4][16] , \REGISTERS[4][15] , \REGISTERS[4][14] ,
         \REGISTERS[4][13] , \REGISTERS[4][12] , \REGISTERS[4][11] ,
         \REGISTERS[4][10] , \REGISTERS[4][9] , \REGISTERS[4][8] ,
         \REGISTERS[4][7] , \REGISTERS[4][6] , \REGISTERS[4][5] ,
         \REGISTERS[4][4] , \REGISTERS[4][3] , \REGISTERS[4][2] ,
         \REGISTERS[4][1] , \REGISTERS[4][0] , \REGISTERS[5][31] ,
         \REGISTERS[5][30] , \REGISTERS[5][29] , \REGISTERS[5][28] ,
         \REGISTERS[5][27] , \REGISTERS[5][26] , \REGISTERS[5][25] ,
         \REGISTERS[5][24] , \REGISTERS[5][23] , \REGISTERS[5][22] ,
         \REGISTERS[5][21] , \REGISTERS[5][20] , \REGISTERS[5][19] ,
         \REGISTERS[5][18] , \REGISTERS[5][17] , \REGISTERS[5][16] ,
         \REGISTERS[5][15] , \REGISTERS[5][14] , \REGISTERS[5][13] ,
         \REGISTERS[5][12] , \REGISTERS[5][11] , \REGISTERS[5][10] ,
         \REGISTERS[5][9] , \REGISTERS[5][8] , \REGISTERS[5][7] ,
         \REGISTERS[5][6] , \REGISTERS[5][5] , \REGISTERS[5][4] ,
         \REGISTERS[5][3] , \REGISTERS[5][2] , \REGISTERS[5][1] ,
         \REGISTERS[5][0] , \REGISTERS[7][31] , \REGISTERS[7][30] ,
         \REGISTERS[7][29] , \REGISTERS[7][28] , \REGISTERS[7][27] ,
         \REGISTERS[7][26] , \REGISTERS[7][25] , \REGISTERS[7][24] ,
         \REGISTERS[7][23] , \REGISTERS[7][22] , \REGISTERS[7][21] ,
         \REGISTERS[7][20] , \REGISTERS[7][19] , \REGISTERS[7][18] ,
         \REGISTERS[7][17] , \REGISTERS[7][16] , \REGISTERS[7][15] ,
         \REGISTERS[7][14] , \REGISTERS[7][13] , \REGISTERS[7][12] ,
         \REGISTERS[7][11] , \REGISTERS[7][10] , \REGISTERS[7][9] ,
         \REGISTERS[7][8] , \REGISTERS[7][7] , \REGISTERS[7][6] ,
         \REGISTERS[7][5] , \REGISTERS[7][4] , \REGISTERS[7][3] ,
         \REGISTERS[7][2] , \REGISTERS[7][1] , \REGISTERS[7][0] ,
         \REGISTERS[8][31] , \REGISTERS[8][30] , \REGISTERS[8][29] ,
         \REGISTERS[8][28] , \REGISTERS[8][27] , \REGISTERS[8][26] ,
         \REGISTERS[8][25] , \REGISTERS[8][24] , \REGISTERS[8][23] ,
         \REGISTERS[8][22] , \REGISTERS[8][21] , \REGISTERS[8][20] ,
         \REGISTERS[8][19] , \REGISTERS[8][18] , \REGISTERS[8][17] ,
         \REGISTERS[8][16] , \REGISTERS[8][15] , \REGISTERS[8][14] ,
         \REGISTERS[8][13] , \REGISTERS[8][12] , \REGISTERS[8][11] ,
         \REGISTERS[8][10] , \REGISTERS[8][9] , \REGISTERS[8][8] ,
         \REGISTERS[8][7] , \REGISTERS[8][6] , \REGISTERS[8][5] ,
         \REGISTERS[8][4] , \REGISTERS[8][3] , \REGISTERS[8][2] ,
         \REGISTERS[8][1] , \REGISTERS[8][0] , \REGISTERS[9][31] ,
         \REGISTERS[9][30] , \REGISTERS[9][29] , \REGISTERS[9][28] ,
         \REGISTERS[9][27] , \REGISTERS[9][26] , \REGISTERS[9][25] ,
         \REGISTERS[9][24] , \REGISTERS[9][23] , \REGISTERS[9][22] ,
         \REGISTERS[9][21] , \REGISTERS[9][20] , \REGISTERS[9][19] ,
         \REGISTERS[9][18] , \REGISTERS[9][17] , \REGISTERS[9][16] ,
         \REGISTERS[9][15] , \REGISTERS[9][14] , \REGISTERS[9][13] ,
         \REGISTERS[9][12] , \REGISTERS[9][11] , \REGISTERS[9][10] ,
         \REGISTERS[9][9] , \REGISTERS[9][8] , \REGISTERS[9][7] ,
         \REGISTERS[9][6] , \REGISTERS[9][5] , \REGISTERS[9][4] ,
         \REGISTERS[9][3] , \REGISTERS[9][2] , \REGISTERS[9][1] ,
         \REGISTERS[9][0] , \REGISTERS[10][31] , \REGISTERS[10][30] ,
         \REGISTERS[10][29] , \REGISTERS[10][28] , \REGISTERS[10][27] ,
         \REGISTERS[10][26] , \REGISTERS[10][25] , \REGISTERS[10][24] ,
         \REGISTERS[10][23] , \REGISTERS[10][22] , \REGISTERS[10][21] ,
         \REGISTERS[10][20] , \REGISTERS[10][19] , \REGISTERS[10][18] ,
         \REGISTERS[10][17] , \REGISTERS[10][16] , \REGISTERS[10][15] ,
         \REGISTERS[10][14] , \REGISTERS[10][13] , \REGISTERS[10][12] ,
         \REGISTERS[10][11] , \REGISTERS[10][10] , \REGISTERS[10][9] ,
         \REGISTERS[10][8] , \REGISTERS[10][7] , \REGISTERS[10][6] ,
         \REGISTERS[10][5] , \REGISTERS[10][4] , \REGISTERS[10][3] ,
         \REGISTERS[10][2] , \REGISTERS[10][1] , \REGISTERS[10][0] ,
         \REGISTERS[11][31] , \REGISTERS[11][30] , \REGISTERS[11][29] ,
         \REGISTERS[11][28] , \REGISTERS[11][27] , \REGISTERS[11][26] ,
         \REGISTERS[11][25] , \REGISTERS[11][24] , \REGISTERS[11][23] ,
         \REGISTERS[11][22] , \REGISTERS[11][21] , \REGISTERS[11][20] ,
         \REGISTERS[11][19] , \REGISTERS[11][18] , \REGISTERS[11][17] ,
         \REGISTERS[11][16] , \REGISTERS[11][15] , \REGISTERS[11][14] ,
         \REGISTERS[11][13] , \REGISTERS[11][12] , \REGISTERS[11][11] ,
         \REGISTERS[11][10] , \REGISTERS[11][9] , \REGISTERS[11][8] ,
         \REGISTERS[11][7] , \REGISTERS[11][6] , \REGISTERS[11][5] ,
         \REGISTERS[11][4] , \REGISTERS[11][3] , \REGISTERS[11][2] ,
         \REGISTERS[11][1] , \REGISTERS[11][0] , \REGISTERS[12][31] ,
         \REGISTERS[12][30] , \REGISTERS[12][29] , \REGISTERS[12][28] ,
         \REGISTERS[12][27] , \REGISTERS[12][26] , \REGISTERS[12][25] ,
         \REGISTERS[12][24] , \REGISTERS[12][23] , \REGISTERS[12][22] ,
         \REGISTERS[12][21] , \REGISTERS[12][20] , \REGISTERS[12][19] ,
         \REGISTERS[12][18] , \REGISTERS[12][17] , \REGISTERS[12][16] ,
         \REGISTERS[12][15] , \REGISTERS[12][14] , \REGISTERS[12][13] ,
         \REGISTERS[12][12] , \REGISTERS[12][11] , \REGISTERS[12][10] ,
         \REGISTERS[12][9] , \REGISTERS[12][8] , \REGISTERS[12][7] ,
         \REGISTERS[12][6] , \REGISTERS[12][5] , \REGISTERS[12][4] ,
         \REGISTERS[12][3] , \REGISTERS[12][2] , \REGISTERS[12][1] ,
         \REGISTERS[12][0] , \REGISTERS[13][31] , \REGISTERS[13][30] ,
         \REGISTERS[13][29] , \REGISTERS[13][28] , \REGISTERS[13][27] ,
         \REGISTERS[13][26] , \REGISTERS[13][25] , \REGISTERS[13][24] ,
         \REGISTERS[13][23] , \REGISTERS[13][22] , \REGISTERS[13][21] ,
         \REGISTERS[13][20] , \REGISTERS[13][19] , \REGISTERS[13][18] ,
         \REGISTERS[13][17] , \REGISTERS[13][16] , \REGISTERS[13][15] ,
         \REGISTERS[13][14] , \REGISTERS[13][13] , \REGISTERS[13][12] ,
         \REGISTERS[13][11] , \REGISTERS[13][10] , \REGISTERS[13][9] ,
         \REGISTERS[13][8] , \REGISTERS[13][7] , \REGISTERS[13][6] ,
         \REGISTERS[13][5] , \REGISTERS[13][4] , \REGISTERS[13][3] ,
         \REGISTERS[13][2] , \REGISTERS[13][1] , \REGISTERS[13][0] ,
         \REGISTERS[14][31] , \REGISTERS[14][30] , \REGISTERS[14][29] ,
         \REGISTERS[14][28] , \REGISTERS[14][27] , \REGISTERS[14][26] ,
         \REGISTERS[14][25] , \REGISTERS[14][24] , \REGISTERS[14][23] ,
         \REGISTERS[14][22] , \REGISTERS[14][21] , \REGISTERS[14][20] ,
         \REGISTERS[14][19] , \REGISTERS[14][18] , \REGISTERS[14][17] ,
         \REGISTERS[14][16] , \REGISTERS[14][15] , \REGISTERS[14][14] ,
         \REGISTERS[14][13] , \REGISTERS[14][12] , \REGISTERS[14][11] ,
         \REGISTERS[14][10] , \REGISTERS[14][9] , \REGISTERS[14][8] ,
         \REGISTERS[14][7] , \REGISTERS[14][6] , \REGISTERS[14][5] ,
         \REGISTERS[14][4] , \REGISTERS[14][3] , \REGISTERS[14][2] ,
         \REGISTERS[14][1] , \REGISTERS[14][0] , \REGISTERS[15][31] ,
         \REGISTERS[15][30] , \REGISTERS[15][29] , \REGISTERS[15][28] ,
         \REGISTERS[15][27] , \REGISTERS[15][26] , \REGISTERS[15][25] ,
         \REGISTERS[15][24] , \REGISTERS[15][23] , \REGISTERS[15][22] ,
         \REGISTERS[15][21] , \REGISTERS[15][20] , \REGISTERS[15][19] ,
         \REGISTERS[15][18] , \REGISTERS[15][17] , \REGISTERS[15][16] ,
         \REGISTERS[15][15] , \REGISTERS[15][14] , \REGISTERS[15][13] ,
         \REGISTERS[15][12] , \REGISTERS[15][11] , \REGISTERS[15][10] ,
         \REGISTERS[15][9] , \REGISTERS[15][8] , \REGISTERS[15][7] ,
         \REGISTERS[15][6] , \REGISTERS[15][5] , \REGISTERS[15][4] ,
         \REGISTERS[15][3] , \REGISTERS[15][2] , \REGISTERS[15][1] ,
         \REGISTERS[15][0] , \REGISTERS[16][31] , \REGISTERS[16][30] ,
         \REGISTERS[16][29] , \REGISTERS[16][28] , \REGISTERS[16][27] ,
         \REGISTERS[16][26] , \REGISTERS[16][25] , \REGISTERS[16][24] ,
         \REGISTERS[16][23] , \REGISTERS[16][22] , \REGISTERS[16][21] ,
         \REGISTERS[16][20] , \REGISTERS[16][19] , \REGISTERS[16][18] ,
         \REGISTERS[16][17] , \REGISTERS[16][16] , \REGISTERS[16][15] ,
         \REGISTERS[16][14] , \REGISTERS[16][13] , \REGISTERS[16][12] ,
         \REGISTERS[16][11] , \REGISTERS[16][10] , \REGISTERS[16][9] ,
         \REGISTERS[16][8] , \REGISTERS[16][7] , \REGISTERS[16][6] ,
         \REGISTERS[16][5] , \REGISTERS[16][4] , \REGISTERS[16][3] ,
         \REGISTERS[16][2] , \REGISTERS[16][1] , \REGISTERS[16][0] ,
         \REGISTERS[17][31] , \REGISTERS[17][30] , \REGISTERS[17][29] ,
         \REGISTERS[17][28] , \REGISTERS[17][27] , \REGISTERS[17][26] ,
         \REGISTERS[17][25] , \REGISTERS[17][24] , \REGISTERS[17][23] ,
         \REGISTERS[17][22] , \REGISTERS[17][21] , \REGISTERS[17][20] ,
         \REGISTERS[17][19] , \REGISTERS[17][18] , \REGISTERS[17][17] ,
         \REGISTERS[17][16] , \REGISTERS[17][15] , \REGISTERS[17][14] ,
         \REGISTERS[17][13] , \REGISTERS[17][12] , \REGISTERS[17][11] ,
         \REGISTERS[17][10] , \REGISTERS[17][9] , \REGISTERS[17][8] ,
         \REGISTERS[17][7] , \REGISTERS[17][6] , \REGISTERS[17][5] ,
         \REGISTERS[17][4] , \REGISTERS[17][3] , \REGISTERS[17][2] ,
         \REGISTERS[17][1] , \REGISTERS[17][0] , \REGISTERS[18][31] ,
         \REGISTERS[18][30] , \REGISTERS[18][29] , \REGISTERS[18][28] ,
         \REGISTERS[18][27] , \REGISTERS[18][26] , \REGISTERS[18][25] ,
         \REGISTERS[18][24] , \REGISTERS[18][23] , \REGISTERS[18][22] ,
         \REGISTERS[18][21] , \REGISTERS[18][20] , \REGISTERS[18][19] ,
         \REGISTERS[18][18] , \REGISTERS[18][17] , \REGISTERS[18][16] ,
         \REGISTERS[18][15] , \REGISTERS[18][14] , \REGISTERS[18][13] ,
         \REGISTERS[18][12] , \REGISTERS[18][11] , \REGISTERS[18][10] ,
         \REGISTERS[18][9] , \REGISTERS[18][8] , \REGISTERS[18][7] ,
         \REGISTERS[18][6] , \REGISTERS[18][5] , \REGISTERS[18][4] ,
         \REGISTERS[18][3] , \REGISTERS[18][2] , \REGISTERS[18][1] ,
         \REGISTERS[18][0] , \REGISTERS[19][31] , \REGISTERS[19][30] ,
         \REGISTERS[19][29] , \REGISTERS[19][28] , \REGISTERS[19][27] ,
         \REGISTERS[19][26] , \REGISTERS[19][25] , \REGISTERS[19][24] ,
         \REGISTERS[19][23] , \REGISTERS[19][22] , \REGISTERS[19][21] ,
         \REGISTERS[19][20] , \REGISTERS[19][19] , \REGISTERS[19][18] ,
         \REGISTERS[19][17] , \REGISTERS[19][16] , \REGISTERS[19][15] ,
         \REGISTERS[19][14] , \REGISTERS[19][13] , \REGISTERS[19][12] ,
         \REGISTERS[19][11] , \REGISTERS[19][10] , \REGISTERS[19][9] ,
         \REGISTERS[19][8] , \REGISTERS[19][7] , \REGISTERS[19][6] ,
         \REGISTERS[19][5] , \REGISTERS[19][4] , \REGISTERS[19][3] ,
         \REGISTERS[19][2] , \REGISTERS[19][1] , \REGISTERS[19][0] ,
         \REGISTERS[20][31] , \REGISTERS[20][30] , \REGISTERS[20][29] ,
         \REGISTERS[20][28] , \REGISTERS[20][27] , \REGISTERS[20][26] ,
         \REGISTERS[20][25] , \REGISTERS[20][24] , \REGISTERS[20][23] ,
         \REGISTERS[20][22] , \REGISTERS[20][21] , \REGISTERS[20][20] ,
         \REGISTERS[20][19] , \REGISTERS[20][18] , \REGISTERS[20][17] ,
         \REGISTERS[20][16] , \REGISTERS[20][15] , \REGISTERS[20][14] ,
         \REGISTERS[20][13] , \REGISTERS[20][12] , \REGISTERS[20][11] ,
         \REGISTERS[20][10] , \REGISTERS[20][9] , \REGISTERS[20][8] ,
         \REGISTERS[20][7] , \REGISTERS[20][6] , \REGISTERS[20][5] ,
         \REGISTERS[20][4] , \REGISTERS[20][3] , \REGISTERS[20][2] ,
         \REGISTERS[20][1] , \REGISTERS[20][0] , \REGISTERS[21][31] ,
         \REGISTERS[21][30] , \REGISTERS[21][29] , \REGISTERS[21][28] ,
         \REGISTERS[21][27] , \REGISTERS[21][26] , \REGISTERS[21][25] ,
         \REGISTERS[21][24] , \REGISTERS[21][23] , \REGISTERS[21][22] ,
         \REGISTERS[21][21] , \REGISTERS[21][20] , \REGISTERS[21][19] ,
         \REGISTERS[21][18] , \REGISTERS[21][17] , \REGISTERS[21][16] ,
         \REGISTERS[21][15] , \REGISTERS[21][14] , \REGISTERS[21][13] ,
         \REGISTERS[21][12] , \REGISTERS[21][11] , \REGISTERS[21][10] ,
         \REGISTERS[21][9] , \REGISTERS[21][8] , \REGISTERS[21][7] ,
         \REGISTERS[21][6] , \REGISTERS[21][5] , \REGISTERS[21][4] ,
         \REGISTERS[21][3] , \REGISTERS[21][2] , \REGISTERS[21][1] ,
         \REGISTERS[21][0] , \REGISTERS[22][31] , \REGISTERS[22][30] ,
         \REGISTERS[22][29] , \REGISTERS[22][28] , \REGISTERS[22][27] ,
         \REGISTERS[22][26] , \REGISTERS[22][25] , \REGISTERS[22][24] ,
         \REGISTERS[22][23] , \REGISTERS[22][22] , \REGISTERS[22][21] ,
         \REGISTERS[22][20] , \REGISTERS[22][19] , \REGISTERS[22][18] ,
         \REGISTERS[22][17] , \REGISTERS[22][16] , \REGISTERS[22][15] ,
         \REGISTERS[22][14] , \REGISTERS[22][13] , \REGISTERS[22][12] ,
         \REGISTERS[22][11] , \REGISTERS[22][10] , \REGISTERS[22][9] ,
         \REGISTERS[22][8] , \REGISTERS[22][7] , \REGISTERS[22][6] ,
         \REGISTERS[22][5] , \REGISTERS[22][4] , \REGISTERS[22][3] ,
         \REGISTERS[22][2] , \REGISTERS[22][1] , \REGISTERS[22][0] ,
         \REGISTERS[23][31] , \REGISTERS[23][30] , \REGISTERS[23][29] ,
         \REGISTERS[23][28] , \REGISTERS[23][27] , \REGISTERS[23][26] ,
         \REGISTERS[23][25] , \REGISTERS[23][24] , \REGISTERS[23][23] ,
         \REGISTERS[23][22] , \REGISTERS[23][21] , \REGISTERS[23][20] ,
         \REGISTERS[23][19] , \REGISTERS[23][18] , \REGISTERS[23][17] ,
         \REGISTERS[23][16] , \REGISTERS[23][15] , \REGISTERS[23][14] ,
         \REGISTERS[23][13] , \REGISTERS[23][12] , \REGISTERS[23][11] ,
         \REGISTERS[23][10] , \REGISTERS[23][9] , \REGISTERS[23][8] ,
         \REGISTERS[23][7] , \REGISTERS[23][6] , \REGISTERS[23][5] ,
         \REGISTERS[23][4] , \REGISTERS[23][3] , \REGISTERS[23][2] ,
         \REGISTERS[23][1] , \REGISTERS[23][0] , \REGISTERS[24][31] ,
         \REGISTERS[24][30] , \REGISTERS[24][29] , \REGISTERS[24][28] ,
         \REGISTERS[24][27] , \REGISTERS[24][26] , \REGISTERS[24][25] ,
         \REGISTERS[24][24] , \REGISTERS[24][23] , \REGISTERS[24][22] ,
         \REGISTERS[24][21] , \REGISTERS[24][20] , \REGISTERS[24][19] ,
         \REGISTERS[24][18] , \REGISTERS[24][17] , \REGISTERS[24][16] ,
         \REGISTERS[24][15] , \REGISTERS[24][14] , \REGISTERS[24][13] ,
         \REGISTERS[24][12] , \REGISTERS[24][11] , \REGISTERS[24][10] ,
         \REGISTERS[24][9] , \REGISTERS[24][8] , \REGISTERS[24][7] ,
         \REGISTERS[24][6] , \REGISTERS[24][5] , \REGISTERS[24][4] ,
         \REGISTERS[24][3] , \REGISTERS[24][2] , \REGISTERS[24][1] ,
         \REGISTERS[24][0] , \REGISTERS[25][31] , \REGISTERS[25][30] ,
         \REGISTERS[25][29] , \REGISTERS[25][28] , \REGISTERS[25][27] ,
         \REGISTERS[25][26] , \REGISTERS[25][25] , \REGISTERS[25][24] ,
         \REGISTERS[25][23] , \REGISTERS[25][22] , \REGISTERS[25][21] ,
         \REGISTERS[25][20] , \REGISTERS[25][19] , \REGISTERS[25][18] ,
         \REGISTERS[25][17] , \REGISTERS[25][16] , \REGISTERS[25][15] ,
         \REGISTERS[25][14] , \REGISTERS[25][13] , \REGISTERS[25][12] ,
         \REGISTERS[25][11] , \REGISTERS[25][10] , \REGISTERS[25][9] ,
         \REGISTERS[25][8] , \REGISTERS[25][7] , \REGISTERS[25][6] ,
         \REGISTERS[25][5] , \REGISTERS[25][4] , \REGISTERS[25][3] ,
         \REGISTERS[25][2] , \REGISTERS[25][1] , \REGISTERS[25][0] ,
         \REGISTERS[26][31] , \REGISTERS[26][30] , \REGISTERS[26][29] ,
         \REGISTERS[26][28] , \REGISTERS[26][27] , \REGISTERS[26][26] ,
         \REGISTERS[26][25] , \REGISTERS[26][24] , \REGISTERS[26][23] ,
         \REGISTERS[26][22] , \REGISTERS[26][21] , \REGISTERS[26][20] ,
         \REGISTERS[26][19] , \REGISTERS[26][18] , \REGISTERS[26][17] ,
         \REGISTERS[26][16] , \REGISTERS[26][15] , \REGISTERS[26][14] ,
         \REGISTERS[26][13] , \REGISTERS[26][12] , \REGISTERS[26][11] ,
         \REGISTERS[26][10] , \REGISTERS[26][9] , \REGISTERS[26][8] ,
         \REGISTERS[26][7] , \REGISTERS[26][6] , \REGISTERS[26][5] ,
         \REGISTERS[26][4] , \REGISTERS[26][3] , \REGISTERS[26][2] ,
         \REGISTERS[26][1] , \REGISTERS[26][0] , \REGISTERS[27][31] ,
         \REGISTERS[27][30] , \REGISTERS[27][29] , \REGISTERS[27][28] ,
         \REGISTERS[27][27] , \REGISTERS[27][26] , \REGISTERS[27][25] ,
         \REGISTERS[27][24] , \REGISTERS[27][23] , \REGISTERS[27][22] ,
         \REGISTERS[27][21] , \REGISTERS[27][20] , \REGISTERS[27][19] ,
         \REGISTERS[27][18] , \REGISTERS[27][17] , \REGISTERS[27][16] ,
         \REGISTERS[27][15] , \REGISTERS[27][14] , \REGISTERS[27][13] ,
         \REGISTERS[27][12] , \REGISTERS[27][11] , \REGISTERS[27][10] ,
         \REGISTERS[27][9] , \REGISTERS[27][8] , \REGISTERS[27][7] ,
         \REGISTERS[27][6] , \REGISTERS[27][5] , \REGISTERS[27][4] ,
         \REGISTERS[27][3] , \REGISTERS[27][2] , \REGISTERS[27][1] ,
         \REGISTERS[27][0] , \REGISTERS[28][31] , \REGISTERS[28][30] ,
         \REGISTERS[28][29] , \REGISTERS[28][28] , \REGISTERS[28][27] ,
         \REGISTERS[28][26] , \REGISTERS[28][25] , \REGISTERS[28][24] ,
         \REGISTERS[28][23] , \REGISTERS[28][22] , \REGISTERS[28][21] ,
         \REGISTERS[28][20] , \REGISTERS[28][19] , \REGISTERS[28][18] ,
         \REGISTERS[28][17] , \REGISTERS[28][16] , \REGISTERS[28][15] ,
         \REGISTERS[28][14] , \REGISTERS[28][13] , \REGISTERS[28][12] ,
         \REGISTERS[28][11] , \REGISTERS[28][10] , \REGISTERS[28][9] ,
         \REGISTERS[28][8] , \REGISTERS[28][7] , \REGISTERS[28][6] ,
         \REGISTERS[28][5] , \REGISTERS[28][4] , \REGISTERS[28][3] ,
         \REGISTERS[28][2] , \REGISTERS[28][1] , \REGISTERS[28][0] ,
         \REGISTERS[29][31] , \REGISTERS[29][30] , \REGISTERS[29][29] ,
         \REGISTERS[29][28] , \REGISTERS[29][27] , \REGISTERS[29][26] ,
         \REGISTERS[29][25] , \REGISTERS[29][24] , \REGISTERS[29][23] ,
         \REGISTERS[29][22] , \REGISTERS[29][21] , \REGISTERS[29][20] ,
         \REGISTERS[29][19] , \REGISTERS[29][18] , \REGISTERS[29][17] ,
         \REGISTERS[29][16] , \REGISTERS[29][15] , \REGISTERS[29][14] ,
         \REGISTERS[29][13] , \REGISTERS[29][12] , \REGISTERS[29][11] ,
         \REGISTERS[29][10] , \REGISTERS[29][9] , \REGISTERS[29][8] ,
         \REGISTERS[29][7] , \REGISTERS[29][6] , \REGISTERS[29][5] ,
         \REGISTERS[29][4] , \REGISTERS[29][3] , \REGISTERS[29][2] ,
         \REGISTERS[29][1] , \REGISTERS[29][0] , \REGISTERS[30][31] ,
         \REGISTERS[30][30] , \REGISTERS[30][29] , \REGISTERS[30][28] ,
         \REGISTERS[30][27] , \REGISTERS[30][26] , \REGISTERS[30][25] ,
         \REGISTERS[30][24] , \REGISTERS[30][23] , \REGISTERS[30][22] ,
         \REGISTERS[30][21] , \REGISTERS[30][20] , \REGISTERS[30][19] ,
         \REGISTERS[30][18] , \REGISTERS[30][17] , \REGISTERS[30][16] ,
         \REGISTERS[30][15] , \REGISTERS[30][14] , \REGISTERS[30][13] ,
         \REGISTERS[30][12] , \REGISTERS[30][11] , \REGISTERS[30][10] ,
         \REGISTERS[30][9] , \REGISTERS[30][8] , \REGISTERS[30][7] ,
         \REGISTERS[30][6] , \REGISTERS[30][5] , \REGISTERS[30][4] ,
         \REGISTERS[30][3] , \REGISTERS[30][2] , \REGISTERS[30][1] ,
         \REGISTERS[30][0] , \REGISTERS[31][31] , \REGISTERS[31][30] ,
         \REGISTERS[31][29] , \REGISTERS[31][28] , \REGISTERS[31][27] ,
         \REGISTERS[31][26] , \REGISTERS[31][25] , \REGISTERS[31][24] ,
         \REGISTERS[31][23] , \REGISTERS[31][22] , \REGISTERS[31][21] ,
         \REGISTERS[31][20] , \REGISTERS[31][19] , \REGISTERS[31][18] ,
         \REGISTERS[31][17] , \REGISTERS[31][16] , \REGISTERS[31][15] ,
         \REGISTERS[31][14] , \REGISTERS[31][13] , \REGISTERS[31][12] ,
         \REGISTERS[31][11] , \REGISTERS[31][10] , \REGISTERS[31][9] ,
         \REGISTERS[31][8] , \REGISTERS[31][7] , \REGISTERS[31][6] ,
         \REGISTERS[31][5] , \REGISTERS[31][4] , \REGISTERS[31][3] ,
         \REGISTERS[31][2] , \REGISTERS[31][1] , \REGISTERS[31][0] , N409,
         N410, N411, N412, N413, N414, N415, N416, N417, N418, N419, N420,
         N421, N422, N423, N424, N425, N426, N427, N428, N429, N430, N431,
         N432, N433, N434, N435, N436, N437, N438, N439, net18859, net18865,
         net18870, net18875, net18880, net18885, net18890, net18895, net18900,
         net18905, net18910, net18915, net18920, net18925, net18930, net18935,
         net18940, net18945, net18950, net18955, net18960, net18965, net18970,
         net18975, net18980, net18985, net18990, net18995, net19000, net19005,
         net19010, n1, n2, n3, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531;

  SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_0 \clk_gate_REGISTERS_reg[1]  ( 
        .CLK(CLK), .EN(N439), .ENCLK(net18859), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_30 \clk_gate_REGISTERS_reg[2]  ( 
        .CLK(CLK), .EN(N438), .ENCLK(net18865), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_29 \clk_gate_REGISTERS_reg[3]  ( 
        .CLK(CLK), .EN(N437), .ENCLK(net18870), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_28 \clk_gate_REGISTERS_reg[4]  ( 
        .CLK(CLK), .EN(N436), .ENCLK(net18875), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_27 \clk_gate_REGISTERS_reg[5]  ( 
        .CLK(CLK), .EN(N435), .ENCLK(net18880), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_26 \clk_gate_REGISTERS_reg[6]  ( 
        .CLK(CLK), .EN(N434), .ENCLK(net18885), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_25 \clk_gate_REGISTERS_reg[7]  ( 
        .CLK(CLK), .EN(N433), .ENCLK(net18890), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_24 \clk_gate_REGISTERS_reg[8]  ( 
        .CLK(CLK), .EN(N432), .ENCLK(net18895), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_23 \clk_gate_REGISTERS_reg[9]  ( 
        .CLK(CLK), .EN(N431), .ENCLK(net18900), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_22 \clk_gate_REGISTERS_reg[10]  ( 
        .CLK(CLK), .EN(N430), .ENCLK(net18905), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_21 \clk_gate_REGISTERS_reg[11]  ( 
        .CLK(CLK), .EN(N429), .ENCLK(net18910), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_20 \clk_gate_REGISTERS_reg[12]  ( 
        .CLK(CLK), .EN(N428), .ENCLK(net18915), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_19 \clk_gate_REGISTERS_reg[13]  ( 
        .CLK(CLK), .EN(N427), .ENCLK(net18920), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_18 \clk_gate_REGISTERS_reg[14]  ( 
        .CLK(CLK), .EN(N426), .ENCLK(net18925), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_17 \clk_gate_REGISTERS_reg[15]  ( 
        .CLK(CLK), .EN(N425), .ENCLK(net18930), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_16 \clk_gate_REGISTERS_reg[16]  ( 
        .CLK(CLK), .EN(N424), .ENCLK(net18935), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_15 \clk_gate_REGISTERS_reg[17]  ( 
        .CLK(CLK), .EN(N423), .ENCLK(net18940), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_14 \clk_gate_REGISTERS_reg[18]  ( 
        .CLK(CLK), .EN(N422), .ENCLK(net18945), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_13 \clk_gate_REGISTERS_reg[19]  ( 
        .CLK(CLK), .EN(N421), .ENCLK(net18950), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_12 \clk_gate_REGISTERS_reg[20]  ( 
        .CLK(CLK), .EN(N420), .ENCLK(net18955), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_11 \clk_gate_REGISTERS_reg[21]  ( 
        .CLK(CLK), .EN(N419), .ENCLK(net18960), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_10 \clk_gate_REGISTERS_reg[22]  ( 
        .CLK(CLK), .EN(N418), .ENCLK(net18965), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_9 \clk_gate_REGISTERS_reg[23]  ( 
        .CLK(CLK), .EN(N417), .ENCLK(net18970), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_8 \clk_gate_REGISTERS_reg[24]  ( 
        .CLK(CLK), .EN(N416), .ENCLK(net18975), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_7 \clk_gate_REGISTERS_reg[25]  ( 
        .CLK(CLK), .EN(N415), .ENCLK(net18980), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_6 \clk_gate_REGISTERS_reg[26]  ( 
        .CLK(CLK), .EN(N414), .ENCLK(net18985), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_5 \clk_gate_REGISTERS_reg[27]  ( 
        .CLK(CLK), .EN(N413), .ENCLK(net18990), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_4 \clk_gate_REGISTERS_reg[28]  ( 
        .CLK(CLK), .EN(N412), .ENCLK(net18995), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_3 \clk_gate_REGISTERS_reg[29]  ( 
        .CLK(CLK), .EN(N411), .ENCLK(net19000), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_2 \clk_gate_REGISTERS_reg[30]  ( 
        .CLK(CLK), .EN(N410), .ENCLK(net19005), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_RF_N_bit32_N_reg32_1 \clk_gate_REGISTERS_reg[31]  ( 
        .CLK(CLK), .EN(N409), .ENCLK(net19010), .TE(1'b0) );
  DFFR_X1 \REGISTERS_reg[1][31]  ( .D(DATA_IN[31]), .CK(net18859), .RN(RST), 
        .Q(\REGISTERS[1][31] ) );
  DFFR_X1 \REGISTERS_reg[1][30]  ( .D(DATA_IN[30]), .CK(net18859), .RN(RST), 
        .Q(\REGISTERS[1][30] ) );
  DFFR_X1 \REGISTERS_reg[1][29]  ( .D(DATA_IN[29]), .CK(net18859), .RN(RST), 
        .Q(\REGISTERS[1][29] ) );
  DFFR_X1 \REGISTERS_reg[1][28]  ( .D(DATA_IN[28]), .CK(net18859), .RN(RST), 
        .Q(\REGISTERS[1][28] ) );
  DFFR_X1 \REGISTERS_reg[1][27]  ( .D(DATA_IN[27]), .CK(net18859), .RN(RST), 
        .Q(\REGISTERS[1][27] ) );
  DFFR_X1 \REGISTERS_reg[1][26]  ( .D(DATA_IN[26]), .CK(net18859), .RN(RST), 
        .Q(\REGISTERS[1][26] ) );
  DFFR_X1 \REGISTERS_reg[1][25]  ( .D(DATA_IN[25]), .CK(net18859), .RN(RST), 
        .Q(\REGISTERS[1][25] ) );
  DFFR_X1 \REGISTERS_reg[1][24]  ( .D(DATA_IN[24]), .CK(net18859), .RN(RST), 
        .Q(\REGISTERS[1][24] ) );
  DFFR_X1 \REGISTERS_reg[1][23]  ( .D(DATA_IN[23]), .CK(net18859), .RN(RST), 
        .Q(\REGISTERS[1][23] ) );
  DFFR_X1 \REGISTERS_reg[1][22]  ( .D(DATA_IN[22]), .CK(net18859), .RN(RST), 
        .Q(\REGISTERS[1][22] ) );
  DFFR_X1 \REGISTERS_reg[1][21]  ( .D(DATA_IN[21]), .CK(net18859), .RN(RST), 
        .Q(\REGISTERS[1][21] ) );
  DFFR_X1 \REGISTERS_reg[1][20]  ( .D(DATA_IN[20]), .CK(net18859), .RN(RST), 
        .Q(\REGISTERS[1][20] ) );
  DFFR_X1 \REGISTERS_reg[1][19]  ( .D(DATA_IN[19]), .CK(net18859), .RN(RST), 
        .Q(\REGISTERS[1][19] ) );
  DFFR_X1 \REGISTERS_reg[1][18]  ( .D(DATA_IN[18]), .CK(net18859), .RN(RST), 
        .Q(\REGISTERS[1][18] ) );
  DFFR_X1 \REGISTERS_reg[1][17]  ( .D(DATA_IN[17]), .CK(net18859), .RN(RST), 
        .Q(\REGISTERS[1][17] ) );
  DFFR_X1 \REGISTERS_reg[1][16]  ( .D(DATA_IN[16]), .CK(net18859), .RN(RST), 
        .Q(\REGISTERS[1][16] ) );
  DFFR_X1 \REGISTERS_reg[1][15]  ( .D(DATA_IN[15]), .CK(net18859), .RN(RST), 
        .Q(\REGISTERS[1][15] ) );
  DFFR_X1 \REGISTERS_reg[1][14]  ( .D(DATA_IN[14]), .CK(net18859), .RN(RST), 
        .Q(\REGISTERS[1][14] ) );
  DFFR_X1 \REGISTERS_reg[1][13]  ( .D(DATA_IN[13]), .CK(net18859), .RN(RST), 
        .Q(\REGISTERS[1][13] ) );
  DFFR_X1 \REGISTERS_reg[1][12]  ( .D(DATA_IN[12]), .CK(net18859), .RN(RST), 
        .Q(\REGISTERS[1][12] ) );
  DFFR_X1 \REGISTERS_reg[1][11]  ( .D(DATA_IN[11]), .CK(net18859), .RN(RST), 
        .Q(\REGISTERS[1][11] ) );
  DFFR_X1 \REGISTERS_reg[1][10]  ( .D(DATA_IN[10]), .CK(net18859), .RN(RST), 
        .Q(\REGISTERS[1][10] ) );
  DFFR_X1 \REGISTERS_reg[1][9]  ( .D(DATA_IN[9]), .CK(net18859), .RN(RST), .Q(
        \REGISTERS[1][9] ) );
  DFFR_X1 \REGISTERS_reg[1][8]  ( .D(DATA_IN[8]), .CK(net18859), .RN(RST), .Q(
        \REGISTERS[1][8] ) );
  DFFR_X1 \REGISTERS_reg[1][7]  ( .D(DATA_IN[7]), .CK(net18859), .RN(RST), .Q(
        \REGISTERS[1][7] ) );
  DFFR_X1 \REGISTERS_reg[1][6]  ( .D(DATA_IN[6]), .CK(net18859), .RN(RST), .Q(
        \REGISTERS[1][6] ) );
  DFFR_X1 \REGISTERS_reg[1][5]  ( .D(DATA_IN[5]), .CK(net18859), .RN(RST), .Q(
        \REGISTERS[1][5] ) );
  DFFR_X1 \REGISTERS_reg[1][4]  ( .D(DATA_IN[4]), .CK(net18859), .RN(RST), .Q(
        \REGISTERS[1][4] ) );
  DFFR_X1 \REGISTERS_reg[1][3]  ( .D(DATA_IN[3]), .CK(net18859), .RN(RST), .Q(
        \REGISTERS[1][3] ) );
  DFFR_X1 \REGISTERS_reg[1][2]  ( .D(DATA_IN[2]), .CK(net18859), .RN(RST), .Q(
        \REGISTERS[1][2] ) );
  DFFR_X1 \REGISTERS_reg[1][1]  ( .D(DATA_IN[1]), .CK(net18859), .RN(RST), .Q(
        \REGISTERS[1][1] ) );
  DFFR_X1 \REGISTERS_reg[1][0]  ( .D(DATA_IN[0]), .CK(net18859), .RN(RST), .Q(
        \REGISTERS[1][0] ) );
  DFFR_X1 \REGISTERS_reg[2][31]  ( .D(DATA_IN[31]), .CK(net18865), .RN(RST), 
        .Q(\REGISTERS[2][31] ) );
  DFFR_X1 \REGISTERS_reg[2][30]  ( .D(DATA_IN[30]), .CK(net18865), .RN(RST), 
        .Q(\REGISTERS[2][30] ) );
  DFFR_X1 \REGISTERS_reg[2][29]  ( .D(DATA_IN[29]), .CK(net18865), .RN(RST), 
        .Q(\REGISTERS[2][29] ) );
  DFFR_X1 \REGISTERS_reg[2][28]  ( .D(DATA_IN[28]), .CK(net18865), .RN(RST), 
        .Q(\REGISTERS[2][28] ) );
  DFFR_X1 \REGISTERS_reg[2][27]  ( .D(DATA_IN[27]), .CK(net18865), .RN(RST), 
        .Q(\REGISTERS[2][27] ) );
  DFFR_X1 \REGISTERS_reg[2][26]  ( .D(DATA_IN[26]), .CK(net18865), .RN(RST), 
        .Q(\REGISTERS[2][26] ) );
  DFFR_X1 \REGISTERS_reg[2][25]  ( .D(DATA_IN[25]), .CK(net18865), .RN(RST), 
        .Q(\REGISTERS[2][25] ) );
  DFFR_X1 \REGISTERS_reg[2][24]  ( .D(DATA_IN[24]), .CK(net18865), .RN(RST), 
        .Q(\REGISTERS[2][24] ) );
  DFFR_X1 \REGISTERS_reg[2][23]  ( .D(DATA_IN[23]), .CK(net18865), .RN(RST), 
        .Q(\REGISTERS[2][23] ) );
  DFFR_X1 \REGISTERS_reg[2][22]  ( .D(DATA_IN[22]), .CK(net18865), .RN(RST), 
        .Q(\REGISTERS[2][22] ) );
  DFFR_X1 \REGISTERS_reg[2][21]  ( .D(DATA_IN[21]), .CK(net18865), .RN(RST), 
        .Q(\REGISTERS[2][21] ) );
  DFFR_X1 \REGISTERS_reg[2][20]  ( .D(DATA_IN[20]), .CK(net18865), .RN(RST), 
        .Q(\REGISTERS[2][20] ) );
  DFFR_X1 \REGISTERS_reg[2][19]  ( .D(DATA_IN[19]), .CK(net18865), .RN(RST), 
        .Q(\REGISTERS[2][19] ) );
  DFFR_X1 \REGISTERS_reg[2][18]  ( .D(DATA_IN[18]), .CK(net18865), .RN(RST), 
        .Q(\REGISTERS[2][18] ) );
  DFFR_X1 \REGISTERS_reg[2][17]  ( .D(DATA_IN[17]), .CK(net18865), .RN(RST), 
        .Q(\REGISTERS[2][17] ) );
  DFFR_X1 \REGISTERS_reg[2][16]  ( .D(DATA_IN[16]), .CK(net18865), .RN(RST), 
        .Q(\REGISTERS[2][16] ) );
  DFFR_X1 \REGISTERS_reg[2][15]  ( .D(DATA_IN[15]), .CK(net18865), .RN(RST), 
        .Q(\REGISTERS[2][15] ) );
  DFFR_X1 \REGISTERS_reg[2][14]  ( .D(DATA_IN[14]), .CK(net18865), .RN(RST), 
        .Q(\REGISTERS[2][14] ) );
  DFFR_X1 \REGISTERS_reg[2][13]  ( .D(DATA_IN[13]), .CK(net18865), .RN(RST), 
        .Q(\REGISTERS[2][13] ) );
  DFFR_X1 \REGISTERS_reg[2][12]  ( .D(DATA_IN[12]), .CK(net18865), .RN(RST), 
        .Q(\REGISTERS[2][12] ) );
  DFFR_X1 \REGISTERS_reg[2][11]  ( .D(DATA_IN[11]), .CK(net18865), .RN(RST), 
        .Q(\REGISTERS[2][11] ) );
  DFFR_X1 \REGISTERS_reg[2][10]  ( .D(DATA_IN[10]), .CK(net18865), .RN(RST), 
        .Q(\REGISTERS[2][10] ) );
  DFFR_X1 \REGISTERS_reg[2][9]  ( .D(DATA_IN[9]), .CK(net18865), .RN(RST), .Q(
        \REGISTERS[2][9] ) );
  DFFR_X1 \REGISTERS_reg[2][8]  ( .D(DATA_IN[8]), .CK(net18865), .RN(RST), .Q(
        \REGISTERS[2][8] ) );
  DFFR_X1 \REGISTERS_reg[2][7]  ( .D(DATA_IN[7]), .CK(net18865), .RN(RST), .Q(
        \REGISTERS[2][7] ) );
  DFFR_X1 \REGISTERS_reg[2][6]  ( .D(DATA_IN[6]), .CK(net18865), .RN(RST), .Q(
        \REGISTERS[2][6] ) );
  DFFR_X1 \REGISTERS_reg[2][5]  ( .D(DATA_IN[5]), .CK(net18865), .RN(RST), .Q(
        \REGISTERS[2][5] ) );
  DFFR_X1 \REGISTERS_reg[2][4]  ( .D(DATA_IN[4]), .CK(net18865), .RN(RST), .Q(
        \REGISTERS[2][4] ) );
  DFFR_X1 \REGISTERS_reg[2][3]  ( .D(DATA_IN[3]), .CK(net18865), .RN(RST), .Q(
        \REGISTERS[2][3] ) );
  DFFR_X1 \REGISTERS_reg[2][2]  ( .D(DATA_IN[2]), .CK(net18865), .RN(RST), .Q(
        \REGISTERS[2][2] ) );
  DFFR_X1 \REGISTERS_reg[2][1]  ( .D(DATA_IN[1]), .CK(net18865), .RN(RST), .Q(
        \REGISTERS[2][1] ) );
  DFFR_X1 \REGISTERS_reg[2][0]  ( .D(DATA_IN[0]), .CK(net18865), .RN(RST), .Q(
        \REGISTERS[2][0] ) );
  DFFR_X1 \REGISTERS_reg[3][31]  ( .D(DATA_IN[31]), .CK(net18870), .RN(RST), 
        .Q(\REGISTERS[3][31] ) );
  DFFR_X1 \REGISTERS_reg[3][30]  ( .D(DATA_IN[30]), .CK(net18870), .RN(RST), 
        .Q(\REGISTERS[3][30] ) );
  DFFR_X1 \REGISTERS_reg[3][29]  ( .D(DATA_IN[29]), .CK(net18870), .RN(RST), 
        .Q(\REGISTERS[3][29] ) );
  DFFR_X1 \REGISTERS_reg[3][28]  ( .D(DATA_IN[28]), .CK(net18870), .RN(RST), 
        .Q(\REGISTERS[3][28] ) );
  DFFR_X1 \REGISTERS_reg[3][27]  ( .D(DATA_IN[27]), .CK(net18870), .RN(RST), 
        .Q(\REGISTERS[3][27] ) );
  DFFR_X1 \REGISTERS_reg[3][26]  ( .D(DATA_IN[26]), .CK(net18870), .RN(RST), 
        .Q(\REGISTERS[3][26] ) );
  DFFR_X1 \REGISTERS_reg[3][25]  ( .D(DATA_IN[25]), .CK(net18870), .RN(RST), 
        .Q(\REGISTERS[3][25] ) );
  DFFR_X1 \REGISTERS_reg[3][24]  ( .D(DATA_IN[24]), .CK(net18870), .RN(RST), 
        .Q(\REGISTERS[3][24] ) );
  DFFR_X1 \REGISTERS_reg[3][23]  ( .D(DATA_IN[23]), .CK(net18870), .RN(RST), 
        .Q(\REGISTERS[3][23] ) );
  DFFR_X1 \REGISTERS_reg[3][22]  ( .D(DATA_IN[22]), .CK(net18870), .RN(RST), 
        .Q(\REGISTERS[3][22] ) );
  DFFR_X1 \REGISTERS_reg[3][21]  ( .D(DATA_IN[21]), .CK(net18870), .RN(RST), 
        .Q(\REGISTERS[3][21] ) );
  DFFR_X1 \REGISTERS_reg[3][20]  ( .D(DATA_IN[20]), .CK(net18870), .RN(RST), 
        .Q(\REGISTERS[3][20] ) );
  DFFR_X1 \REGISTERS_reg[3][19]  ( .D(DATA_IN[19]), .CK(net18870), .RN(RST), 
        .Q(\REGISTERS[3][19] ) );
  DFFR_X1 \REGISTERS_reg[3][18]  ( .D(DATA_IN[18]), .CK(net18870), .RN(RST), 
        .Q(\REGISTERS[3][18] ) );
  DFFR_X1 \REGISTERS_reg[3][17]  ( .D(DATA_IN[17]), .CK(net18870), .RN(RST), 
        .Q(\REGISTERS[3][17] ) );
  DFFR_X1 \REGISTERS_reg[3][16]  ( .D(DATA_IN[16]), .CK(net18870), .RN(RST), 
        .Q(\REGISTERS[3][16] ) );
  DFFR_X1 \REGISTERS_reg[3][15]  ( .D(DATA_IN[15]), .CK(net18870), .RN(RST), 
        .Q(\REGISTERS[3][15] ) );
  DFFR_X1 \REGISTERS_reg[3][14]  ( .D(DATA_IN[14]), .CK(net18870), .RN(RST), 
        .Q(\REGISTERS[3][14] ) );
  DFFR_X1 \REGISTERS_reg[3][13]  ( .D(DATA_IN[13]), .CK(net18870), .RN(RST), 
        .Q(\REGISTERS[3][13] ) );
  DFFR_X1 \REGISTERS_reg[3][12]  ( .D(DATA_IN[12]), .CK(net18870), .RN(RST), 
        .Q(\REGISTERS[3][12] ) );
  DFFR_X1 \REGISTERS_reg[3][11]  ( .D(DATA_IN[11]), .CK(net18870), .RN(RST), 
        .Q(\REGISTERS[3][11] ) );
  DFFR_X1 \REGISTERS_reg[3][10]  ( .D(DATA_IN[10]), .CK(net18870), .RN(RST), 
        .Q(\REGISTERS[3][10] ) );
  DFFR_X1 \REGISTERS_reg[3][9]  ( .D(DATA_IN[9]), .CK(net18870), .RN(RST), .Q(
        \REGISTERS[3][9] ) );
  DFFR_X1 \REGISTERS_reg[3][8]  ( .D(DATA_IN[8]), .CK(net18870), .RN(RST), .Q(
        \REGISTERS[3][8] ) );
  DFFR_X1 \REGISTERS_reg[3][7]  ( .D(DATA_IN[7]), .CK(net18870), .RN(RST), .Q(
        \REGISTERS[3][7] ) );
  DFFR_X1 \REGISTERS_reg[3][6]  ( .D(DATA_IN[6]), .CK(net18870), .RN(RST), .Q(
        \REGISTERS[3][6] ) );
  DFFR_X1 \REGISTERS_reg[3][5]  ( .D(DATA_IN[5]), .CK(net18870), .RN(RST), .Q(
        \REGISTERS[3][5] ) );
  DFFR_X1 \REGISTERS_reg[3][4]  ( .D(DATA_IN[4]), .CK(net18870), .RN(RST), .Q(
        \REGISTERS[3][4] ) );
  DFFR_X1 \REGISTERS_reg[3][3]  ( .D(DATA_IN[3]), .CK(net18870), .RN(RST), .Q(
        \REGISTERS[3][3] ) );
  DFFR_X1 \REGISTERS_reg[3][2]  ( .D(DATA_IN[2]), .CK(net18870), .RN(RST), .Q(
        \REGISTERS[3][2] ) );
  DFFR_X1 \REGISTERS_reg[3][1]  ( .D(DATA_IN[1]), .CK(net18870), .RN(RST), .Q(
        \REGISTERS[3][1] ) );
  DFFR_X1 \REGISTERS_reg[3][0]  ( .D(DATA_IN[0]), .CK(net18870), .RN(RST), .Q(
        \REGISTERS[3][0] ) );
  DFFR_X1 \REGISTERS_reg[4][31]  ( .D(DATA_IN[31]), .CK(net18875), .RN(RST), 
        .Q(\REGISTERS[4][31] ) );
  DFFR_X1 \REGISTERS_reg[4][30]  ( .D(DATA_IN[30]), .CK(net18875), .RN(RST), 
        .Q(\REGISTERS[4][30] ) );
  DFFR_X1 \REGISTERS_reg[4][29]  ( .D(DATA_IN[29]), .CK(net18875), .RN(RST), 
        .Q(\REGISTERS[4][29] ) );
  DFFR_X1 \REGISTERS_reg[4][28]  ( .D(DATA_IN[28]), .CK(net18875), .RN(RST), 
        .Q(\REGISTERS[4][28] ) );
  DFFR_X1 \REGISTERS_reg[4][27]  ( .D(DATA_IN[27]), .CK(net18875), .RN(RST), 
        .Q(\REGISTERS[4][27] ) );
  DFFR_X1 \REGISTERS_reg[4][26]  ( .D(DATA_IN[26]), .CK(net18875), .RN(RST), 
        .Q(\REGISTERS[4][26] ) );
  DFFR_X1 \REGISTERS_reg[4][25]  ( .D(DATA_IN[25]), .CK(net18875), .RN(RST), 
        .Q(\REGISTERS[4][25] ) );
  DFFR_X1 \REGISTERS_reg[4][24]  ( .D(DATA_IN[24]), .CK(net18875), .RN(RST), 
        .Q(\REGISTERS[4][24] ) );
  DFFR_X1 \REGISTERS_reg[4][23]  ( .D(DATA_IN[23]), .CK(net18875), .RN(RST), 
        .Q(\REGISTERS[4][23] ) );
  DFFR_X1 \REGISTERS_reg[4][22]  ( .D(DATA_IN[22]), .CK(net18875), .RN(RST), 
        .Q(\REGISTERS[4][22] ) );
  DFFR_X1 \REGISTERS_reg[4][21]  ( .D(DATA_IN[21]), .CK(net18875), .RN(RST), 
        .Q(\REGISTERS[4][21] ) );
  DFFR_X1 \REGISTERS_reg[4][20]  ( .D(DATA_IN[20]), .CK(net18875), .RN(RST), 
        .Q(\REGISTERS[4][20] ) );
  DFFR_X1 \REGISTERS_reg[4][19]  ( .D(DATA_IN[19]), .CK(net18875), .RN(RST), 
        .Q(\REGISTERS[4][19] ) );
  DFFR_X1 \REGISTERS_reg[4][18]  ( .D(DATA_IN[18]), .CK(net18875), .RN(RST), 
        .Q(\REGISTERS[4][18] ) );
  DFFR_X1 \REGISTERS_reg[4][17]  ( .D(DATA_IN[17]), .CK(net18875), .RN(RST), 
        .Q(\REGISTERS[4][17] ) );
  DFFR_X1 \REGISTERS_reg[4][16]  ( .D(DATA_IN[16]), .CK(net18875), .RN(RST), 
        .Q(\REGISTERS[4][16] ) );
  DFFR_X1 \REGISTERS_reg[4][15]  ( .D(DATA_IN[15]), .CK(net18875), .RN(RST), 
        .Q(\REGISTERS[4][15] ) );
  DFFR_X1 \REGISTERS_reg[4][14]  ( .D(DATA_IN[14]), .CK(net18875), .RN(RST), 
        .Q(\REGISTERS[4][14] ) );
  DFFR_X1 \REGISTERS_reg[4][13]  ( .D(DATA_IN[13]), .CK(net18875), .RN(RST), 
        .Q(\REGISTERS[4][13] ) );
  DFFR_X1 \REGISTERS_reg[4][12]  ( .D(DATA_IN[12]), .CK(net18875), .RN(RST), 
        .Q(\REGISTERS[4][12] ) );
  DFFR_X1 \REGISTERS_reg[4][11]  ( .D(DATA_IN[11]), .CK(net18875), .RN(RST), 
        .Q(\REGISTERS[4][11] ) );
  DFFR_X1 \REGISTERS_reg[4][10]  ( .D(DATA_IN[10]), .CK(net18875), .RN(RST), 
        .Q(\REGISTERS[4][10] ) );
  DFFR_X1 \REGISTERS_reg[4][9]  ( .D(DATA_IN[9]), .CK(net18875), .RN(RST), .Q(
        \REGISTERS[4][9] ) );
  DFFR_X1 \REGISTERS_reg[4][8]  ( .D(DATA_IN[8]), .CK(net18875), .RN(RST), .Q(
        \REGISTERS[4][8] ) );
  DFFR_X1 \REGISTERS_reg[4][7]  ( .D(DATA_IN[7]), .CK(net18875), .RN(RST), .Q(
        \REGISTERS[4][7] ) );
  DFFR_X1 \REGISTERS_reg[4][6]  ( .D(DATA_IN[6]), .CK(net18875), .RN(RST), .Q(
        \REGISTERS[4][6] ) );
  DFFR_X1 \REGISTERS_reg[4][5]  ( .D(DATA_IN[5]), .CK(net18875), .RN(RST), .Q(
        \REGISTERS[4][5] ) );
  DFFR_X1 \REGISTERS_reg[4][4]  ( .D(DATA_IN[4]), .CK(net18875), .RN(RST), .Q(
        \REGISTERS[4][4] ) );
  DFFR_X1 \REGISTERS_reg[4][3]  ( .D(DATA_IN[3]), .CK(net18875), .RN(RST), .Q(
        \REGISTERS[4][3] ) );
  DFFR_X1 \REGISTERS_reg[4][2]  ( .D(DATA_IN[2]), .CK(net18875), .RN(RST), .Q(
        \REGISTERS[4][2] ) );
  DFFR_X1 \REGISTERS_reg[4][1]  ( .D(DATA_IN[1]), .CK(net18875), .RN(RST), .Q(
        \REGISTERS[4][1] ) );
  DFFR_X1 \REGISTERS_reg[4][0]  ( .D(DATA_IN[0]), .CK(net18875), .RN(RST), .Q(
        \REGISTERS[4][0] ) );
  DFFR_X1 \REGISTERS_reg[5][31]  ( .D(DATA_IN[31]), .CK(net18880), .RN(RST), 
        .Q(\REGISTERS[5][31] ) );
  DFFR_X1 \REGISTERS_reg[5][30]  ( .D(DATA_IN[30]), .CK(net18880), .RN(RST), 
        .Q(\REGISTERS[5][30] ) );
  DFFR_X1 \REGISTERS_reg[5][29]  ( .D(DATA_IN[29]), .CK(net18880), .RN(RST), 
        .Q(\REGISTERS[5][29] ) );
  DFFR_X1 \REGISTERS_reg[5][28]  ( .D(DATA_IN[28]), .CK(net18880), .RN(RST), 
        .Q(\REGISTERS[5][28] ) );
  DFFR_X1 \REGISTERS_reg[5][27]  ( .D(DATA_IN[27]), .CK(net18880), .RN(RST), 
        .Q(\REGISTERS[5][27] ) );
  DFFR_X1 \REGISTERS_reg[5][26]  ( .D(DATA_IN[26]), .CK(net18880), .RN(RST), 
        .Q(\REGISTERS[5][26] ) );
  DFFR_X1 \REGISTERS_reg[5][25]  ( .D(DATA_IN[25]), .CK(net18880), .RN(RST), 
        .Q(\REGISTERS[5][25] ) );
  DFFR_X1 \REGISTERS_reg[5][24]  ( .D(DATA_IN[24]), .CK(net18880), .RN(RST), 
        .Q(\REGISTERS[5][24] ) );
  DFFR_X1 \REGISTERS_reg[5][23]  ( .D(DATA_IN[23]), .CK(net18880), .RN(RST), 
        .Q(\REGISTERS[5][23] ) );
  DFFR_X1 \REGISTERS_reg[5][22]  ( .D(DATA_IN[22]), .CK(net18880), .RN(RST), 
        .Q(\REGISTERS[5][22] ) );
  DFFR_X1 \REGISTERS_reg[5][21]  ( .D(DATA_IN[21]), .CK(net18880), .RN(RST), 
        .Q(\REGISTERS[5][21] ) );
  DFFR_X1 \REGISTERS_reg[5][20]  ( .D(DATA_IN[20]), .CK(net18880), .RN(RST), 
        .Q(\REGISTERS[5][20] ) );
  DFFR_X1 \REGISTERS_reg[5][19]  ( .D(DATA_IN[19]), .CK(net18880), .RN(RST), 
        .Q(\REGISTERS[5][19] ) );
  DFFR_X1 \REGISTERS_reg[5][18]  ( .D(DATA_IN[18]), .CK(net18880), .RN(RST), 
        .Q(\REGISTERS[5][18] ) );
  DFFR_X1 \REGISTERS_reg[5][17]  ( .D(DATA_IN[17]), .CK(net18880), .RN(RST), 
        .Q(\REGISTERS[5][17] ) );
  DFFR_X1 \REGISTERS_reg[5][16]  ( .D(DATA_IN[16]), .CK(net18880), .RN(RST), 
        .Q(\REGISTERS[5][16] ) );
  DFFR_X1 \REGISTERS_reg[5][15]  ( .D(DATA_IN[15]), .CK(net18880), .RN(RST), 
        .Q(\REGISTERS[5][15] ) );
  DFFR_X1 \REGISTERS_reg[5][14]  ( .D(DATA_IN[14]), .CK(net18880), .RN(RST), 
        .Q(\REGISTERS[5][14] ) );
  DFFR_X1 \REGISTERS_reg[5][13]  ( .D(DATA_IN[13]), .CK(net18880), .RN(RST), 
        .Q(\REGISTERS[5][13] ) );
  DFFR_X1 \REGISTERS_reg[5][12]  ( .D(DATA_IN[12]), .CK(net18880), .RN(RST), 
        .Q(\REGISTERS[5][12] ) );
  DFFR_X1 \REGISTERS_reg[5][11]  ( .D(DATA_IN[11]), .CK(net18880), .RN(RST), 
        .Q(\REGISTERS[5][11] ) );
  DFFR_X1 \REGISTERS_reg[5][10]  ( .D(DATA_IN[10]), .CK(net18880), .RN(RST), 
        .Q(\REGISTERS[5][10] ) );
  DFFR_X1 \REGISTERS_reg[5][9]  ( .D(DATA_IN[9]), .CK(net18880), .RN(RST), .Q(
        \REGISTERS[5][9] ) );
  DFFR_X1 \REGISTERS_reg[5][8]  ( .D(DATA_IN[8]), .CK(net18880), .RN(RST), .Q(
        \REGISTERS[5][8] ) );
  DFFR_X1 \REGISTERS_reg[5][7]  ( .D(DATA_IN[7]), .CK(net18880), .RN(RST), .Q(
        \REGISTERS[5][7] ) );
  DFFR_X1 \REGISTERS_reg[5][6]  ( .D(DATA_IN[6]), .CK(net18880), .RN(RST), .Q(
        \REGISTERS[5][6] ) );
  DFFR_X1 \REGISTERS_reg[5][5]  ( .D(DATA_IN[5]), .CK(net18880), .RN(RST), .Q(
        \REGISTERS[5][5] ) );
  DFFR_X1 \REGISTERS_reg[5][4]  ( .D(DATA_IN[4]), .CK(net18880), .RN(RST), .Q(
        \REGISTERS[5][4] ) );
  DFFR_X1 \REGISTERS_reg[5][3]  ( .D(DATA_IN[3]), .CK(net18880), .RN(RST), .Q(
        \REGISTERS[5][3] ) );
  DFFR_X1 \REGISTERS_reg[5][2]  ( .D(DATA_IN[2]), .CK(net18880), .RN(RST), .Q(
        \REGISTERS[5][2] ) );
  DFFR_X1 \REGISTERS_reg[5][1]  ( .D(DATA_IN[1]), .CK(net18880), .RN(RST), .Q(
        \REGISTERS[5][1] ) );
  DFFR_X1 \REGISTERS_reg[5][0]  ( .D(DATA_IN[0]), .CK(net18880), .RN(RST), .Q(
        \REGISTERS[5][0] ) );
  DFFR_X1 \REGISTERS_reg[6][31]  ( .D(DATA_IN[31]), .CK(net18885), .RN(RST), 
        .QN(n62) );
  DFFR_X1 \REGISTERS_reg[6][30]  ( .D(DATA_IN[30]), .CK(net18885), .RN(RST), 
        .QN(n61) );
  DFFR_X1 \REGISTERS_reg[6][29]  ( .D(DATA_IN[29]), .CK(net18885), .RN(RST), 
        .QN(n59) );
  DFFR_X1 \REGISTERS_reg[6][28]  ( .D(DATA_IN[28]), .CK(net18885), .RN(RST), 
        .QN(n58) );
  DFFR_X1 \REGISTERS_reg[6][27]  ( .D(DATA_IN[27]), .CK(net18885), .RN(RST), 
        .QN(n57) );
  DFFR_X1 \REGISTERS_reg[6][26]  ( .D(DATA_IN[26]), .CK(net18885), .RN(RST), 
        .QN(n56) );
  DFFR_X1 \REGISTERS_reg[6][25]  ( .D(DATA_IN[25]), .CK(net18885), .RN(RST), 
        .QN(n55) );
  DFFR_X1 \REGISTERS_reg[6][24]  ( .D(DATA_IN[24]), .CK(net18885), .RN(RST), 
        .QN(n54) );
  DFFR_X1 \REGISTERS_reg[6][23]  ( .D(DATA_IN[23]), .CK(net18885), .RN(RST), 
        .QN(n53) );
  DFFR_X1 \REGISTERS_reg[6][22]  ( .D(DATA_IN[22]), .CK(net18885), .RN(RST), 
        .QN(n52) );
  DFFR_X1 \REGISTERS_reg[6][21]  ( .D(DATA_IN[21]), .CK(net18885), .RN(RST), 
        .QN(n51) );
  DFFR_X1 \REGISTERS_reg[6][20]  ( .D(DATA_IN[20]), .CK(net18885), .RN(RST), 
        .QN(n50) );
  DFFR_X1 \REGISTERS_reg[6][19]  ( .D(DATA_IN[19]), .CK(net18885), .RN(RST), 
        .QN(n48) );
  DFFR_X1 \REGISTERS_reg[6][18]  ( .D(DATA_IN[18]), .CK(net18885), .RN(RST), 
        .QN(n47) );
  DFFR_X1 \REGISTERS_reg[6][17]  ( .D(DATA_IN[17]), .CK(net18885), .RN(RST), 
        .QN(n46) );
  DFFR_X1 \REGISTERS_reg[6][16]  ( .D(DATA_IN[16]), .CK(net18885), .RN(RST), 
        .QN(n45) );
  DFFR_X1 \REGISTERS_reg[6][15]  ( .D(DATA_IN[15]), .CK(net18885), .RN(RST), 
        .QN(n44) );
  DFFR_X1 \REGISTERS_reg[6][14]  ( .D(DATA_IN[14]), .CK(net18885), .RN(RST), 
        .QN(n43) );
  DFFR_X1 \REGISTERS_reg[6][13]  ( .D(DATA_IN[13]), .CK(net18885), .RN(RST), 
        .QN(n42) );
  DFFR_X1 \REGISTERS_reg[6][12]  ( .D(DATA_IN[12]), .CK(net18885), .RN(RST), 
        .QN(n41) );
  DFFR_X1 \REGISTERS_reg[6][11]  ( .D(DATA_IN[11]), .CK(net18885), .RN(RST), 
        .QN(n40) );
  DFFR_X1 \REGISTERS_reg[6][10]  ( .D(DATA_IN[10]), .CK(net18885), .RN(RST), 
        .QN(n39) );
  DFFR_X1 \REGISTERS_reg[6][9]  ( .D(DATA_IN[9]), .CK(net18885), .RN(RST), 
        .QN(n69) );
  DFFR_X1 \REGISTERS_reg[6][8]  ( .D(DATA_IN[8]), .CK(net18885), .RN(RST), 
        .QN(n68) );
  DFFR_X1 \REGISTERS_reg[6][7]  ( .D(DATA_IN[7]), .CK(net18885), .RN(RST), 
        .QN(n67) );
  DFFR_X1 \REGISTERS_reg[6][6]  ( .D(DATA_IN[6]), .CK(net18885), .RN(RST), 
        .QN(n66) );
  DFFR_X1 \REGISTERS_reg[6][5]  ( .D(DATA_IN[5]), .CK(net18885), .RN(RST), 
        .QN(n65) );
  DFFR_X1 \REGISTERS_reg[6][4]  ( .D(DATA_IN[4]), .CK(net18885), .RN(RST), 
        .QN(n64) );
  DFFR_X1 \REGISTERS_reg[6][3]  ( .D(DATA_IN[3]), .CK(net18885), .RN(RST), 
        .QN(n63) );
  DFFR_X1 \REGISTERS_reg[6][2]  ( .D(DATA_IN[2]), .CK(net18885), .RN(RST), 
        .QN(n60) );
  DFFR_X1 \REGISTERS_reg[6][1]  ( .D(DATA_IN[1]), .CK(net18885), .RN(RST), 
        .QN(n49) );
  DFFR_X1 \REGISTERS_reg[6][0]  ( .D(DATA_IN[0]), .CK(net18885), .RN(RST), 
        .QN(n38) );
  DFFR_X1 \REGISTERS_reg[7][31]  ( .D(DATA_IN[31]), .CK(net18890), .RN(RST), 
        .Q(\REGISTERS[7][31] ) );
  DFFR_X1 \REGISTERS_reg[7][30]  ( .D(DATA_IN[30]), .CK(net18890), .RN(RST), 
        .Q(\REGISTERS[7][30] ) );
  DFFR_X1 \REGISTERS_reg[7][29]  ( .D(DATA_IN[29]), .CK(net18890), .RN(RST), 
        .Q(\REGISTERS[7][29] ) );
  DFFR_X1 \REGISTERS_reg[7][28]  ( .D(DATA_IN[28]), .CK(net18890), .RN(RST), 
        .Q(\REGISTERS[7][28] ) );
  DFFR_X1 \REGISTERS_reg[7][27]  ( .D(DATA_IN[27]), .CK(net18890), .RN(RST), 
        .Q(\REGISTERS[7][27] ) );
  DFFR_X1 \REGISTERS_reg[7][26]  ( .D(DATA_IN[26]), .CK(net18890), .RN(RST), 
        .Q(\REGISTERS[7][26] ) );
  DFFR_X1 \REGISTERS_reg[7][25]  ( .D(DATA_IN[25]), .CK(net18890), .RN(RST), 
        .Q(\REGISTERS[7][25] ) );
  DFFR_X1 \REGISTERS_reg[7][24]  ( .D(DATA_IN[24]), .CK(net18890), .RN(RST), 
        .Q(\REGISTERS[7][24] ) );
  DFFR_X1 \REGISTERS_reg[7][23]  ( .D(DATA_IN[23]), .CK(net18890), .RN(RST), 
        .Q(\REGISTERS[7][23] ) );
  DFFR_X1 \REGISTERS_reg[7][22]  ( .D(DATA_IN[22]), .CK(net18890), .RN(RST), 
        .Q(\REGISTERS[7][22] ) );
  DFFR_X1 \REGISTERS_reg[7][21]  ( .D(DATA_IN[21]), .CK(net18890), .RN(RST), 
        .Q(\REGISTERS[7][21] ) );
  DFFR_X1 \REGISTERS_reg[7][20]  ( .D(DATA_IN[20]), .CK(net18890), .RN(RST), 
        .Q(\REGISTERS[7][20] ) );
  DFFR_X1 \REGISTERS_reg[7][19]  ( .D(DATA_IN[19]), .CK(net18890), .RN(RST), 
        .Q(\REGISTERS[7][19] ) );
  DFFR_X1 \REGISTERS_reg[7][18]  ( .D(DATA_IN[18]), .CK(net18890), .RN(RST), 
        .Q(\REGISTERS[7][18] ) );
  DFFR_X1 \REGISTERS_reg[7][17]  ( .D(DATA_IN[17]), .CK(net18890), .RN(RST), 
        .Q(\REGISTERS[7][17] ) );
  DFFR_X1 \REGISTERS_reg[7][16]  ( .D(DATA_IN[16]), .CK(net18890), .RN(RST), 
        .Q(\REGISTERS[7][16] ) );
  DFFR_X1 \REGISTERS_reg[7][15]  ( .D(DATA_IN[15]), .CK(net18890), .RN(RST), 
        .Q(\REGISTERS[7][15] ) );
  DFFR_X1 \REGISTERS_reg[7][14]  ( .D(DATA_IN[14]), .CK(net18890), .RN(RST), 
        .Q(\REGISTERS[7][14] ) );
  DFFR_X1 \REGISTERS_reg[7][13]  ( .D(DATA_IN[13]), .CK(net18890), .RN(RST), 
        .Q(\REGISTERS[7][13] ) );
  DFFR_X1 \REGISTERS_reg[7][12]  ( .D(DATA_IN[12]), .CK(net18890), .RN(RST), 
        .Q(\REGISTERS[7][12] ) );
  DFFR_X1 \REGISTERS_reg[7][11]  ( .D(DATA_IN[11]), .CK(net18890), .RN(RST), 
        .Q(\REGISTERS[7][11] ) );
  DFFR_X1 \REGISTERS_reg[7][10]  ( .D(DATA_IN[10]), .CK(net18890), .RN(RST), 
        .Q(\REGISTERS[7][10] ) );
  DFFR_X1 \REGISTERS_reg[7][9]  ( .D(DATA_IN[9]), .CK(net18890), .RN(RST), .Q(
        \REGISTERS[7][9] ) );
  DFFR_X1 \REGISTERS_reg[7][8]  ( .D(DATA_IN[8]), .CK(net18890), .RN(RST), .Q(
        \REGISTERS[7][8] ) );
  DFFR_X1 \REGISTERS_reg[7][7]  ( .D(DATA_IN[7]), .CK(net18890), .RN(RST), .Q(
        \REGISTERS[7][7] ) );
  DFFR_X1 \REGISTERS_reg[7][6]  ( .D(DATA_IN[6]), .CK(net18890), .RN(RST), .Q(
        \REGISTERS[7][6] ) );
  DFFR_X1 \REGISTERS_reg[7][5]  ( .D(DATA_IN[5]), .CK(net18890), .RN(RST), .Q(
        \REGISTERS[7][5] ) );
  DFFR_X1 \REGISTERS_reg[7][4]  ( .D(DATA_IN[4]), .CK(net18890), .RN(RST), .Q(
        \REGISTERS[7][4] ) );
  DFFR_X1 \REGISTERS_reg[7][3]  ( .D(DATA_IN[3]), .CK(net18890), .RN(RST), .Q(
        \REGISTERS[7][3] ) );
  DFFR_X1 \REGISTERS_reg[7][2]  ( .D(DATA_IN[2]), .CK(net18890), .RN(RST), .Q(
        \REGISTERS[7][2] ) );
  DFFR_X1 \REGISTERS_reg[7][1]  ( .D(DATA_IN[1]), .CK(net18890), .RN(RST), .Q(
        \REGISTERS[7][1] ) );
  DFFR_X1 \REGISTERS_reg[7][0]  ( .D(DATA_IN[0]), .CK(net18890), .RN(RST), .Q(
        \REGISTERS[7][0] ) );
  DFFR_X1 \REGISTERS_reg[8][31]  ( .D(DATA_IN[31]), .CK(net18895), .RN(RST), 
        .Q(\REGISTERS[8][31] ) );
  DFFR_X1 \REGISTERS_reg[8][30]  ( .D(DATA_IN[30]), .CK(net18895), .RN(RST), 
        .Q(\REGISTERS[8][30] ) );
  DFFR_X1 \REGISTERS_reg[8][29]  ( .D(DATA_IN[29]), .CK(net18895), .RN(RST), 
        .Q(\REGISTERS[8][29] ) );
  DFFR_X1 \REGISTERS_reg[8][28]  ( .D(DATA_IN[28]), .CK(net18895), .RN(RST), 
        .Q(\REGISTERS[8][28] ) );
  DFFR_X1 \REGISTERS_reg[8][27]  ( .D(DATA_IN[27]), .CK(net18895), .RN(RST), 
        .Q(\REGISTERS[8][27] ) );
  DFFR_X1 \REGISTERS_reg[8][26]  ( .D(DATA_IN[26]), .CK(net18895), .RN(RST), 
        .Q(\REGISTERS[8][26] ) );
  DFFR_X1 \REGISTERS_reg[8][25]  ( .D(DATA_IN[25]), .CK(net18895), .RN(RST), 
        .Q(\REGISTERS[8][25] ) );
  DFFR_X1 \REGISTERS_reg[8][24]  ( .D(DATA_IN[24]), .CK(net18895), .RN(RST), 
        .Q(\REGISTERS[8][24] ) );
  DFFR_X1 \REGISTERS_reg[8][23]  ( .D(DATA_IN[23]), .CK(net18895), .RN(RST), 
        .Q(\REGISTERS[8][23] ) );
  DFFR_X1 \REGISTERS_reg[8][22]  ( .D(DATA_IN[22]), .CK(net18895), .RN(RST), 
        .Q(\REGISTERS[8][22] ) );
  DFFR_X1 \REGISTERS_reg[8][21]  ( .D(DATA_IN[21]), .CK(net18895), .RN(RST), 
        .Q(\REGISTERS[8][21] ) );
  DFFR_X1 \REGISTERS_reg[8][20]  ( .D(DATA_IN[20]), .CK(net18895), .RN(RST), 
        .Q(\REGISTERS[8][20] ) );
  DFFR_X1 \REGISTERS_reg[8][19]  ( .D(DATA_IN[19]), .CK(net18895), .RN(RST), 
        .Q(\REGISTERS[8][19] ) );
  DFFR_X1 \REGISTERS_reg[8][18]  ( .D(DATA_IN[18]), .CK(net18895), .RN(RST), 
        .Q(\REGISTERS[8][18] ) );
  DFFR_X1 \REGISTERS_reg[8][17]  ( .D(DATA_IN[17]), .CK(net18895), .RN(RST), 
        .Q(\REGISTERS[8][17] ) );
  DFFR_X1 \REGISTERS_reg[8][16]  ( .D(DATA_IN[16]), .CK(net18895), .RN(RST), 
        .Q(\REGISTERS[8][16] ) );
  DFFR_X1 \REGISTERS_reg[8][15]  ( .D(DATA_IN[15]), .CK(net18895), .RN(RST), 
        .Q(\REGISTERS[8][15] ) );
  DFFR_X1 \REGISTERS_reg[8][14]  ( .D(DATA_IN[14]), .CK(net18895), .RN(RST), 
        .Q(\REGISTERS[8][14] ) );
  DFFR_X1 \REGISTERS_reg[8][13]  ( .D(DATA_IN[13]), .CK(net18895), .RN(RST), 
        .Q(\REGISTERS[8][13] ) );
  DFFR_X1 \REGISTERS_reg[8][12]  ( .D(DATA_IN[12]), .CK(net18895), .RN(RST), 
        .Q(\REGISTERS[8][12] ) );
  DFFR_X1 \REGISTERS_reg[8][11]  ( .D(DATA_IN[11]), .CK(net18895), .RN(RST), 
        .Q(\REGISTERS[8][11] ) );
  DFFR_X1 \REGISTERS_reg[8][10]  ( .D(DATA_IN[10]), .CK(net18895), .RN(RST), 
        .Q(\REGISTERS[8][10] ) );
  DFFR_X1 \REGISTERS_reg[8][9]  ( .D(DATA_IN[9]), .CK(net18895), .RN(RST), .Q(
        \REGISTERS[8][9] ) );
  DFFR_X1 \REGISTERS_reg[8][8]  ( .D(DATA_IN[8]), .CK(net18895), .RN(RST), .Q(
        \REGISTERS[8][8] ) );
  DFFR_X1 \REGISTERS_reg[8][7]  ( .D(DATA_IN[7]), .CK(net18895), .RN(RST), .Q(
        \REGISTERS[8][7] ) );
  DFFR_X1 \REGISTERS_reg[8][6]  ( .D(DATA_IN[6]), .CK(net18895), .RN(RST), .Q(
        \REGISTERS[8][6] ) );
  DFFR_X1 \REGISTERS_reg[8][5]  ( .D(DATA_IN[5]), .CK(net18895), .RN(RST), .Q(
        \REGISTERS[8][5] ) );
  DFFR_X1 \REGISTERS_reg[8][4]  ( .D(DATA_IN[4]), .CK(net18895), .RN(RST), .Q(
        \REGISTERS[8][4] ) );
  DFFR_X1 \REGISTERS_reg[8][3]  ( .D(DATA_IN[3]), .CK(net18895), .RN(RST), .Q(
        \REGISTERS[8][3] ) );
  DFFR_X1 \REGISTERS_reg[8][2]  ( .D(DATA_IN[2]), .CK(net18895), .RN(RST), .Q(
        \REGISTERS[8][2] ) );
  DFFR_X1 \REGISTERS_reg[8][1]  ( .D(DATA_IN[1]), .CK(net18895), .RN(RST), .Q(
        \REGISTERS[8][1] ) );
  DFFR_X1 \REGISTERS_reg[8][0]  ( .D(DATA_IN[0]), .CK(net18895), .RN(RST), .Q(
        \REGISTERS[8][0] ) );
  DFFR_X1 \REGISTERS_reg[9][31]  ( .D(DATA_IN[31]), .CK(net18900), .RN(RST), 
        .Q(\REGISTERS[9][31] ) );
  DFFR_X1 \REGISTERS_reg[9][30]  ( .D(DATA_IN[30]), .CK(net18900), .RN(RST), 
        .Q(\REGISTERS[9][30] ) );
  DFFR_X1 \REGISTERS_reg[9][29]  ( .D(DATA_IN[29]), .CK(net18900), .RN(RST), 
        .Q(\REGISTERS[9][29] ) );
  DFFR_X1 \REGISTERS_reg[9][28]  ( .D(DATA_IN[28]), .CK(net18900), .RN(RST), 
        .Q(\REGISTERS[9][28] ) );
  DFFR_X1 \REGISTERS_reg[9][27]  ( .D(DATA_IN[27]), .CK(net18900), .RN(RST), 
        .Q(\REGISTERS[9][27] ) );
  DFFR_X1 \REGISTERS_reg[9][26]  ( .D(DATA_IN[26]), .CK(net18900), .RN(RST), 
        .Q(\REGISTERS[9][26] ) );
  DFFR_X1 \REGISTERS_reg[9][25]  ( .D(DATA_IN[25]), .CK(net18900), .RN(RST), 
        .Q(\REGISTERS[9][25] ) );
  DFFR_X1 \REGISTERS_reg[9][24]  ( .D(DATA_IN[24]), .CK(net18900), .RN(RST), 
        .Q(\REGISTERS[9][24] ) );
  DFFR_X1 \REGISTERS_reg[9][23]  ( .D(DATA_IN[23]), .CK(net18900), .RN(RST), 
        .Q(\REGISTERS[9][23] ) );
  DFFR_X1 \REGISTERS_reg[9][22]  ( .D(DATA_IN[22]), .CK(net18900), .RN(RST), 
        .Q(\REGISTERS[9][22] ) );
  DFFR_X1 \REGISTERS_reg[9][21]  ( .D(DATA_IN[21]), .CK(net18900), .RN(RST), 
        .Q(\REGISTERS[9][21] ) );
  DFFR_X1 \REGISTERS_reg[9][20]  ( .D(DATA_IN[20]), .CK(net18900), .RN(RST), 
        .Q(\REGISTERS[9][20] ) );
  DFFR_X1 \REGISTERS_reg[9][19]  ( .D(DATA_IN[19]), .CK(net18900), .RN(RST), 
        .Q(\REGISTERS[9][19] ) );
  DFFR_X1 \REGISTERS_reg[9][18]  ( .D(DATA_IN[18]), .CK(net18900), .RN(RST), 
        .Q(\REGISTERS[9][18] ) );
  DFFR_X1 \REGISTERS_reg[9][17]  ( .D(DATA_IN[17]), .CK(net18900), .RN(RST), 
        .Q(\REGISTERS[9][17] ) );
  DFFR_X1 \REGISTERS_reg[9][16]  ( .D(DATA_IN[16]), .CK(net18900), .RN(RST), 
        .Q(\REGISTERS[9][16] ) );
  DFFR_X1 \REGISTERS_reg[9][15]  ( .D(DATA_IN[15]), .CK(net18900), .RN(RST), 
        .Q(\REGISTERS[9][15] ) );
  DFFR_X1 \REGISTERS_reg[9][14]  ( .D(DATA_IN[14]), .CK(net18900), .RN(RST), 
        .Q(\REGISTERS[9][14] ) );
  DFFR_X1 \REGISTERS_reg[9][13]  ( .D(DATA_IN[13]), .CK(net18900), .RN(RST), 
        .Q(\REGISTERS[9][13] ) );
  DFFR_X1 \REGISTERS_reg[9][12]  ( .D(DATA_IN[12]), .CK(net18900), .RN(RST), 
        .Q(\REGISTERS[9][12] ) );
  DFFR_X1 \REGISTERS_reg[9][11]  ( .D(DATA_IN[11]), .CK(net18900), .RN(RST), 
        .Q(\REGISTERS[9][11] ) );
  DFFR_X1 \REGISTERS_reg[9][10]  ( .D(DATA_IN[10]), .CK(net18900), .RN(RST), 
        .Q(\REGISTERS[9][10] ) );
  DFFR_X1 \REGISTERS_reg[9][9]  ( .D(DATA_IN[9]), .CK(net18900), .RN(RST), .Q(
        \REGISTERS[9][9] ) );
  DFFR_X1 \REGISTERS_reg[9][8]  ( .D(DATA_IN[8]), .CK(net18900), .RN(RST), .Q(
        \REGISTERS[9][8] ) );
  DFFR_X1 \REGISTERS_reg[9][7]  ( .D(DATA_IN[7]), .CK(net18900), .RN(RST), .Q(
        \REGISTERS[9][7] ) );
  DFFR_X1 \REGISTERS_reg[9][6]  ( .D(DATA_IN[6]), .CK(net18900), .RN(RST), .Q(
        \REGISTERS[9][6] ) );
  DFFR_X1 \REGISTERS_reg[9][5]  ( .D(DATA_IN[5]), .CK(net18900), .RN(RST), .Q(
        \REGISTERS[9][5] ) );
  DFFR_X1 \REGISTERS_reg[9][4]  ( .D(DATA_IN[4]), .CK(net18900), .RN(RST), .Q(
        \REGISTERS[9][4] ) );
  DFFR_X1 \REGISTERS_reg[9][3]  ( .D(DATA_IN[3]), .CK(net18900), .RN(RST), .Q(
        \REGISTERS[9][3] ) );
  DFFR_X1 \REGISTERS_reg[9][2]  ( .D(DATA_IN[2]), .CK(net18900), .RN(RST), .Q(
        \REGISTERS[9][2] ) );
  DFFR_X1 \REGISTERS_reg[9][1]  ( .D(DATA_IN[1]), .CK(net18900), .RN(RST), .Q(
        \REGISTERS[9][1] ) );
  DFFR_X1 \REGISTERS_reg[9][0]  ( .D(DATA_IN[0]), .CK(net18900), .RN(RST), .Q(
        \REGISTERS[9][0] ) );
  DFFR_X1 \REGISTERS_reg[10][31]  ( .D(DATA_IN[31]), .CK(net18905), .RN(RST), 
        .Q(\REGISTERS[10][31] ) );
  DFFR_X1 \REGISTERS_reg[10][30]  ( .D(DATA_IN[30]), .CK(net18905), .RN(RST), 
        .Q(\REGISTERS[10][30] ) );
  DFFR_X1 \REGISTERS_reg[10][29]  ( .D(DATA_IN[29]), .CK(net18905), .RN(RST), 
        .Q(\REGISTERS[10][29] ) );
  DFFR_X1 \REGISTERS_reg[10][28]  ( .D(DATA_IN[28]), .CK(net18905), .RN(RST), 
        .Q(\REGISTERS[10][28] ) );
  DFFR_X1 \REGISTERS_reg[10][27]  ( .D(DATA_IN[27]), .CK(net18905), .RN(RST), 
        .Q(\REGISTERS[10][27] ) );
  DFFR_X1 \REGISTERS_reg[10][26]  ( .D(DATA_IN[26]), .CK(net18905), .RN(RST), 
        .Q(\REGISTERS[10][26] ) );
  DFFR_X1 \REGISTERS_reg[10][25]  ( .D(DATA_IN[25]), .CK(net18905), .RN(RST), 
        .Q(\REGISTERS[10][25] ) );
  DFFR_X1 \REGISTERS_reg[10][24]  ( .D(DATA_IN[24]), .CK(net18905), .RN(RST), 
        .Q(\REGISTERS[10][24] ) );
  DFFR_X1 \REGISTERS_reg[10][23]  ( .D(DATA_IN[23]), .CK(net18905), .RN(RST), 
        .Q(\REGISTERS[10][23] ) );
  DFFR_X1 \REGISTERS_reg[10][22]  ( .D(DATA_IN[22]), .CK(net18905), .RN(RST), 
        .Q(\REGISTERS[10][22] ) );
  DFFR_X1 \REGISTERS_reg[10][21]  ( .D(DATA_IN[21]), .CK(net18905), .RN(RST), 
        .Q(\REGISTERS[10][21] ) );
  DFFR_X1 \REGISTERS_reg[10][20]  ( .D(DATA_IN[20]), .CK(net18905), .RN(RST), 
        .Q(\REGISTERS[10][20] ) );
  DFFR_X1 \REGISTERS_reg[10][19]  ( .D(DATA_IN[19]), .CK(net18905), .RN(RST), 
        .Q(\REGISTERS[10][19] ) );
  DFFR_X1 \REGISTERS_reg[10][18]  ( .D(DATA_IN[18]), .CK(net18905), .RN(RST), 
        .Q(\REGISTERS[10][18] ) );
  DFFR_X1 \REGISTERS_reg[10][17]  ( .D(DATA_IN[17]), .CK(net18905), .RN(RST), 
        .Q(\REGISTERS[10][17] ) );
  DFFR_X1 \REGISTERS_reg[10][16]  ( .D(DATA_IN[16]), .CK(net18905), .RN(RST), 
        .Q(\REGISTERS[10][16] ) );
  DFFR_X1 \REGISTERS_reg[10][15]  ( .D(DATA_IN[15]), .CK(net18905), .RN(RST), 
        .Q(\REGISTERS[10][15] ) );
  DFFR_X1 \REGISTERS_reg[10][14]  ( .D(DATA_IN[14]), .CK(net18905), .RN(RST), 
        .Q(\REGISTERS[10][14] ) );
  DFFR_X1 \REGISTERS_reg[10][13]  ( .D(DATA_IN[13]), .CK(net18905), .RN(RST), 
        .Q(\REGISTERS[10][13] ) );
  DFFR_X1 \REGISTERS_reg[10][12]  ( .D(DATA_IN[12]), .CK(net18905), .RN(RST), 
        .Q(\REGISTERS[10][12] ) );
  DFFR_X1 \REGISTERS_reg[10][11]  ( .D(DATA_IN[11]), .CK(net18905), .RN(RST), 
        .Q(\REGISTERS[10][11] ) );
  DFFR_X1 \REGISTERS_reg[10][10]  ( .D(DATA_IN[10]), .CK(net18905), .RN(RST), 
        .Q(\REGISTERS[10][10] ) );
  DFFR_X1 \REGISTERS_reg[10][9]  ( .D(DATA_IN[9]), .CK(net18905), .RN(RST), 
        .Q(\REGISTERS[10][9] ) );
  DFFR_X1 \REGISTERS_reg[10][8]  ( .D(DATA_IN[8]), .CK(net18905), .RN(RST), 
        .Q(\REGISTERS[10][8] ) );
  DFFR_X1 \REGISTERS_reg[10][7]  ( .D(DATA_IN[7]), .CK(net18905), .RN(RST), 
        .Q(\REGISTERS[10][7] ) );
  DFFR_X1 \REGISTERS_reg[10][6]  ( .D(DATA_IN[6]), .CK(net18905), .RN(RST), 
        .Q(\REGISTERS[10][6] ) );
  DFFR_X1 \REGISTERS_reg[10][5]  ( .D(DATA_IN[5]), .CK(net18905), .RN(RST), 
        .Q(\REGISTERS[10][5] ) );
  DFFR_X1 \REGISTERS_reg[10][4]  ( .D(DATA_IN[4]), .CK(net18905), .RN(RST), 
        .Q(\REGISTERS[10][4] ) );
  DFFR_X1 \REGISTERS_reg[10][3]  ( .D(DATA_IN[3]), .CK(net18905), .RN(RST), 
        .Q(\REGISTERS[10][3] ) );
  DFFR_X1 \REGISTERS_reg[10][2]  ( .D(DATA_IN[2]), .CK(net18905), .RN(RST), 
        .Q(\REGISTERS[10][2] ) );
  DFFR_X1 \REGISTERS_reg[10][1]  ( .D(DATA_IN[1]), .CK(net18905), .RN(RST), 
        .Q(\REGISTERS[10][1] ) );
  DFFR_X1 \REGISTERS_reg[10][0]  ( .D(DATA_IN[0]), .CK(net18905), .RN(RST), 
        .Q(\REGISTERS[10][0] ) );
  DFFR_X1 \REGISTERS_reg[11][31]  ( .D(DATA_IN[31]), .CK(net18910), .RN(RST), 
        .Q(\REGISTERS[11][31] ) );
  DFFR_X1 \REGISTERS_reg[11][30]  ( .D(DATA_IN[30]), .CK(net18910), .RN(RST), 
        .Q(\REGISTERS[11][30] ) );
  DFFR_X1 \REGISTERS_reg[11][29]  ( .D(DATA_IN[29]), .CK(net18910), .RN(RST), 
        .Q(\REGISTERS[11][29] ) );
  DFFR_X1 \REGISTERS_reg[11][28]  ( .D(DATA_IN[28]), .CK(net18910), .RN(RST), 
        .Q(\REGISTERS[11][28] ) );
  DFFR_X1 \REGISTERS_reg[11][27]  ( .D(DATA_IN[27]), .CK(net18910), .RN(RST), 
        .Q(\REGISTERS[11][27] ) );
  DFFR_X1 \REGISTERS_reg[11][26]  ( .D(DATA_IN[26]), .CK(net18910), .RN(RST), 
        .Q(\REGISTERS[11][26] ) );
  DFFR_X1 \REGISTERS_reg[11][25]  ( .D(DATA_IN[25]), .CK(net18910), .RN(RST), 
        .Q(\REGISTERS[11][25] ) );
  DFFR_X1 \REGISTERS_reg[11][24]  ( .D(DATA_IN[24]), .CK(net18910), .RN(RST), 
        .Q(\REGISTERS[11][24] ) );
  DFFR_X1 \REGISTERS_reg[11][23]  ( .D(DATA_IN[23]), .CK(net18910), .RN(RST), 
        .Q(\REGISTERS[11][23] ) );
  DFFR_X1 \REGISTERS_reg[11][22]  ( .D(DATA_IN[22]), .CK(net18910), .RN(RST), 
        .Q(\REGISTERS[11][22] ) );
  DFFR_X1 \REGISTERS_reg[11][21]  ( .D(DATA_IN[21]), .CK(net18910), .RN(RST), 
        .Q(\REGISTERS[11][21] ) );
  DFFR_X1 \REGISTERS_reg[11][20]  ( .D(DATA_IN[20]), .CK(net18910), .RN(RST), 
        .Q(\REGISTERS[11][20] ) );
  DFFR_X1 \REGISTERS_reg[11][19]  ( .D(DATA_IN[19]), .CK(net18910), .RN(RST), 
        .Q(\REGISTERS[11][19] ) );
  DFFR_X1 \REGISTERS_reg[11][18]  ( .D(DATA_IN[18]), .CK(net18910), .RN(RST), 
        .Q(\REGISTERS[11][18] ) );
  DFFR_X1 \REGISTERS_reg[11][17]  ( .D(DATA_IN[17]), .CK(net18910), .RN(RST), 
        .Q(\REGISTERS[11][17] ) );
  DFFR_X1 \REGISTERS_reg[11][16]  ( .D(DATA_IN[16]), .CK(net18910), .RN(RST), 
        .Q(\REGISTERS[11][16] ) );
  DFFR_X1 \REGISTERS_reg[11][15]  ( .D(DATA_IN[15]), .CK(net18910), .RN(RST), 
        .Q(\REGISTERS[11][15] ) );
  DFFR_X1 \REGISTERS_reg[11][14]  ( .D(DATA_IN[14]), .CK(net18910), .RN(RST), 
        .Q(\REGISTERS[11][14] ) );
  DFFR_X1 \REGISTERS_reg[11][13]  ( .D(DATA_IN[13]), .CK(net18910), .RN(RST), 
        .Q(\REGISTERS[11][13] ) );
  DFFR_X1 \REGISTERS_reg[11][12]  ( .D(DATA_IN[12]), .CK(net18910), .RN(RST), 
        .Q(\REGISTERS[11][12] ) );
  DFFR_X1 \REGISTERS_reg[11][11]  ( .D(DATA_IN[11]), .CK(net18910), .RN(RST), 
        .Q(\REGISTERS[11][11] ) );
  DFFR_X1 \REGISTERS_reg[11][10]  ( .D(DATA_IN[10]), .CK(net18910), .RN(RST), 
        .Q(\REGISTERS[11][10] ) );
  DFFR_X1 \REGISTERS_reg[11][9]  ( .D(DATA_IN[9]), .CK(net18910), .RN(RST), 
        .Q(\REGISTERS[11][9] ) );
  DFFR_X1 \REGISTERS_reg[11][8]  ( .D(DATA_IN[8]), .CK(net18910), .RN(RST), 
        .Q(\REGISTERS[11][8] ) );
  DFFR_X1 \REGISTERS_reg[11][7]  ( .D(DATA_IN[7]), .CK(net18910), .RN(RST), 
        .Q(\REGISTERS[11][7] ) );
  DFFR_X1 \REGISTERS_reg[11][6]  ( .D(DATA_IN[6]), .CK(net18910), .RN(RST), 
        .Q(\REGISTERS[11][6] ) );
  DFFR_X1 \REGISTERS_reg[11][5]  ( .D(DATA_IN[5]), .CK(net18910), .RN(RST), 
        .Q(\REGISTERS[11][5] ) );
  DFFR_X1 \REGISTERS_reg[11][4]  ( .D(DATA_IN[4]), .CK(net18910), .RN(RST), 
        .Q(\REGISTERS[11][4] ) );
  DFFR_X1 \REGISTERS_reg[11][3]  ( .D(DATA_IN[3]), .CK(net18910), .RN(RST), 
        .Q(\REGISTERS[11][3] ) );
  DFFR_X1 \REGISTERS_reg[11][2]  ( .D(DATA_IN[2]), .CK(net18910), .RN(RST), 
        .Q(\REGISTERS[11][2] ) );
  DFFR_X1 \REGISTERS_reg[11][1]  ( .D(DATA_IN[1]), .CK(net18910), .RN(RST), 
        .Q(\REGISTERS[11][1] ) );
  DFFR_X1 \REGISTERS_reg[11][0]  ( .D(DATA_IN[0]), .CK(net18910), .RN(RST), 
        .Q(\REGISTERS[11][0] ) );
  DFFR_X1 \REGISTERS_reg[12][31]  ( .D(DATA_IN[31]), .CK(net18915), .RN(RST), 
        .Q(\REGISTERS[12][31] ) );
  DFFR_X1 \REGISTERS_reg[12][30]  ( .D(DATA_IN[30]), .CK(net18915), .RN(RST), 
        .Q(\REGISTERS[12][30] ) );
  DFFR_X1 \REGISTERS_reg[12][29]  ( .D(DATA_IN[29]), .CK(net18915), .RN(RST), 
        .Q(\REGISTERS[12][29] ) );
  DFFR_X1 \REGISTERS_reg[12][28]  ( .D(DATA_IN[28]), .CK(net18915), .RN(RST), 
        .Q(\REGISTERS[12][28] ) );
  DFFR_X1 \REGISTERS_reg[12][27]  ( .D(DATA_IN[27]), .CK(net18915), .RN(RST), 
        .Q(\REGISTERS[12][27] ) );
  DFFR_X1 \REGISTERS_reg[12][26]  ( .D(DATA_IN[26]), .CK(net18915), .RN(RST), 
        .Q(\REGISTERS[12][26] ) );
  DFFR_X1 \REGISTERS_reg[12][25]  ( .D(DATA_IN[25]), .CK(net18915), .RN(RST), 
        .Q(\REGISTERS[12][25] ) );
  DFFR_X1 \REGISTERS_reg[12][24]  ( .D(DATA_IN[24]), .CK(net18915), .RN(RST), 
        .Q(\REGISTERS[12][24] ) );
  DFFR_X1 \REGISTERS_reg[12][23]  ( .D(DATA_IN[23]), .CK(net18915), .RN(RST), 
        .Q(\REGISTERS[12][23] ) );
  DFFR_X1 \REGISTERS_reg[12][22]  ( .D(DATA_IN[22]), .CK(net18915), .RN(RST), 
        .Q(\REGISTERS[12][22] ) );
  DFFR_X1 \REGISTERS_reg[12][21]  ( .D(DATA_IN[21]), .CK(net18915), .RN(RST), 
        .Q(\REGISTERS[12][21] ) );
  DFFR_X1 \REGISTERS_reg[12][20]  ( .D(DATA_IN[20]), .CK(net18915), .RN(RST), 
        .Q(\REGISTERS[12][20] ) );
  DFFR_X1 \REGISTERS_reg[12][19]  ( .D(DATA_IN[19]), .CK(net18915), .RN(RST), 
        .Q(\REGISTERS[12][19] ) );
  DFFR_X1 \REGISTERS_reg[12][18]  ( .D(DATA_IN[18]), .CK(net18915), .RN(RST), 
        .Q(\REGISTERS[12][18] ) );
  DFFR_X1 \REGISTERS_reg[12][17]  ( .D(DATA_IN[17]), .CK(net18915), .RN(RST), 
        .Q(\REGISTERS[12][17] ) );
  DFFR_X1 \REGISTERS_reg[12][16]  ( .D(DATA_IN[16]), .CK(net18915), .RN(RST), 
        .Q(\REGISTERS[12][16] ) );
  DFFR_X1 \REGISTERS_reg[12][15]  ( .D(DATA_IN[15]), .CK(net18915), .RN(RST), 
        .Q(\REGISTERS[12][15] ) );
  DFFR_X1 \REGISTERS_reg[12][14]  ( .D(DATA_IN[14]), .CK(net18915), .RN(RST), 
        .Q(\REGISTERS[12][14] ) );
  DFFR_X1 \REGISTERS_reg[12][13]  ( .D(DATA_IN[13]), .CK(net18915), .RN(RST), 
        .Q(\REGISTERS[12][13] ) );
  DFFR_X1 \REGISTERS_reg[12][12]  ( .D(DATA_IN[12]), .CK(net18915), .RN(RST), 
        .Q(\REGISTERS[12][12] ) );
  DFFR_X1 \REGISTERS_reg[12][11]  ( .D(DATA_IN[11]), .CK(net18915), .RN(RST), 
        .Q(\REGISTERS[12][11] ) );
  DFFR_X1 \REGISTERS_reg[12][10]  ( .D(DATA_IN[10]), .CK(net18915), .RN(RST), 
        .Q(\REGISTERS[12][10] ) );
  DFFR_X1 \REGISTERS_reg[12][9]  ( .D(DATA_IN[9]), .CK(net18915), .RN(RST), 
        .Q(\REGISTERS[12][9] ) );
  DFFR_X1 \REGISTERS_reg[12][8]  ( .D(DATA_IN[8]), .CK(net18915), .RN(RST), 
        .Q(\REGISTERS[12][8] ) );
  DFFR_X1 \REGISTERS_reg[12][7]  ( .D(DATA_IN[7]), .CK(net18915), .RN(RST), 
        .Q(\REGISTERS[12][7] ) );
  DFFR_X1 \REGISTERS_reg[12][6]  ( .D(DATA_IN[6]), .CK(net18915), .RN(RST), 
        .Q(\REGISTERS[12][6] ) );
  DFFR_X1 \REGISTERS_reg[12][5]  ( .D(DATA_IN[5]), .CK(net18915), .RN(RST), 
        .Q(\REGISTERS[12][5] ) );
  DFFR_X1 \REGISTERS_reg[12][4]  ( .D(DATA_IN[4]), .CK(net18915), .RN(RST), 
        .Q(\REGISTERS[12][4] ) );
  DFFR_X1 \REGISTERS_reg[12][3]  ( .D(DATA_IN[3]), .CK(net18915), .RN(RST), 
        .Q(\REGISTERS[12][3] ) );
  DFFR_X1 \REGISTERS_reg[12][2]  ( .D(DATA_IN[2]), .CK(net18915), .RN(RST), 
        .Q(\REGISTERS[12][2] ) );
  DFFR_X1 \REGISTERS_reg[12][1]  ( .D(DATA_IN[1]), .CK(net18915), .RN(RST), 
        .Q(\REGISTERS[12][1] ) );
  DFFR_X1 \REGISTERS_reg[12][0]  ( .D(DATA_IN[0]), .CK(net18915), .RN(RST), 
        .Q(\REGISTERS[12][0] ) );
  DFFR_X1 \REGISTERS_reg[13][31]  ( .D(DATA_IN[31]), .CK(net18920), .RN(RST), 
        .Q(\REGISTERS[13][31] ) );
  DFFR_X1 \REGISTERS_reg[13][30]  ( .D(DATA_IN[30]), .CK(net18920), .RN(RST), 
        .Q(\REGISTERS[13][30] ) );
  DFFR_X1 \REGISTERS_reg[13][29]  ( .D(DATA_IN[29]), .CK(net18920), .RN(RST), 
        .Q(\REGISTERS[13][29] ) );
  DFFR_X1 \REGISTERS_reg[13][28]  ( .D(DATA_IN[28]), .CK(net18920), .RN(RST), 
        .Q(\REGISTERS[13][28] ) );
  DFFR_X1 \REGISTERS_reg[13][27]  ( .D(DATA_IN[27]), .CK(net18920), .RN(RST), 
        .Q(\REGISTERS[13][27] ) );
  DFFR_X1 \REGISTERS_reg[13][26]  ( .D(DATA_IN[26]), .CK(net18920), .RN(RST), 
        .Q(\REGISTERS[13][26] ) );
  DFFR_X1 \REGISTERS_reg[13][25]  ( .D(DATA_IN[25]), .CK(net18920), .RN(RST), 
        .Q(\REGISTERS[13][25] ) );
  DFFR_X1 \REGISTERS_reg[13][24]  ( .D(DATA_IN[24]), .CK(net18920), .RN(RST), 
        .Q(\REGISTERS[13][24] ) );
  DFFR_X1 \REGISTERS_reg[13][23]  ( .D(DATA_IN[23]), .CK(net18920), .RN(RST), 
        .Q(\REGISTERS[13][23] ) );
  DFFR_X1 \REGISTERS_reg[13][22]  ( .D(DATA_IN[22]), .CK(net18920), .RN(RST), 
        .Q(\REGISTERS[13][22] ) );
  DFFR_X1 \REGISTERS_reg[13][21]  ( .D(DATA_IN[21]), .CK(net18920), .RN(RST), 
        .Q(\REGISTERS[13][21] ) );
  DFFR_X1 \REGISTERS_reg[13][20]  ( .D(DATA_IN[20]), .CK(net18920), .RN(RST), 
        .Q(\REGISTERS[13][20] ) );
  DFFR_X1 \REGISTERS_reg[13][19]  ( .D(DATA_IN[19]), .CK(net18920), .RN(RST), 
        .Q(\REGISTERS[13][19] ) );
  DFFR_X1 \REGISTERS_reg[13][18]  ( .D(DATA_IN[18]), .CK(net18920), .RN(RST), 
        .Q(\REGISTERS[13][18] ) );
  DFFR_X1 \REGISTERS_reg[13][17]  ( .D(DATA_IN[17]), .CK(net18920), .RN(RST), 
        .Q(\REGISTERS[13][17] ) );
  DFFR_X1 \REGISTERS_reg[13][16]  ( .D(DATA_IN[16]), .CK(net18920), .RN(RST), 
        .Q(\REGISTERS[13][16] ) );
  DFFR_X1 \REGISTERS_reg[13][15]  ( .D(DATA_IN[15]), .CK(net18920), .RN(RST), 
        .Q(\REGISTERS[13][15] ) );
  DFFR_X1 \REGISTERS_reg[13][14]  ( .D(DATA_IN[14]), .CK(net18920), .RN(RST), 
        .Q(\REGISTERS[13][14] ) );
  DFFR_X1 \REGISTERS_reg[13][13]  ( .D(DATA_IN[13]), .CK(net18920), .RN(RST), 
        .Q(\REGISTERS[13][13] ) );
  DFFR_X1 \REGISTERS_reg[13][12]  ( .D(DATA_IN[12]), .CK(net18920), .RN(RST), 
        .Q(\REGISTERS[13][12] ) );
  DFFR_X1 \REGISTERS_reg[13][11]  ( .D(DATA_IN[11]), .CK(net18920), .RN(RST), 
        .Q(\REGISTERS[13][11] ) );
  DFFR_X1 \REGISTERS_reg[13][10]  ( .D(DATA_IN[10]), .CK(net18920), .RN(RST), 
        .Q(\REGISTERS[13][10] ) );
  DFFR_X1 \REGISTERS_reg[13][9]  ( .D(DATA_IN[9]), .CK(net18920), .RN(RST), 
        .Q(\REGISTERS[13][9] ) );
  DFFR_X1 \REGISTERS_reg[13][8]  ( .D(DATA_IN[8]), .CK(net18920), .RN(RST), 
        .Q(\REGISTERS[13][8] ) );
  DFFR_X1 \REGISTERS_reg[13][7]  ( .D(DATA_IN[7]), .CK(net18920), .RN(RST), 
        .Q(\REGISTERS[13][7] ) );
  DFFR_X1 \REGISTERS_reg[13][6]  ( .D(DATA_IN[6]), .CK(net18920), .RN(RST), 
        .Q(\REGISTERS[13][6] ) );
  DFFR_X1 \REGISTERS_reg[13][5]  ( .D(DATA_IN[5]), .CK(net18920), .RN(RST), 
        .Q(\REGISTERS[13][5] ) );
  DFFR_X1 \REGISTERS_reg[13][4]  ( .D(DATA_IN[4]), .CK(net18920), .RN(RST), 
        .Q(\REGISTERS[13][4] ) );
  DFFR_X1 \REGISTERS_reg[13][3]  ( .D(DATA_IN[3]), .CK(net18920), .RN(RST), 
        .Q(\REGISTERS[13][3] ) );
  DFFR_X1 \REGISTERS_reg[13][2]  ( .D(DATA_IN[2]), .CK(net18920), .RN(RST), 
        .Q(\REGISTERS[13][2] ) );
  DFFR_X1 \REGISTERS_reg[13][1]  ( .D(DATA_IN[1]), .CK(net18920), .RN(RST), 
        .Q(\REGISTERS[13][1] ) );
  DFFR_X1 \REGISTERS_reg[13][0]  ( .D(DATA_IN[0]), .CK(net18920), .RN(RST), 
        .Q(\REGISTERS[13][0] ) );
  DFFR_X1 \REGISTERS_reg[14][31]  ( .D(DATA_IN[31]), .CK(net18925), .RN(RST), 
        .Q(\REGISTERS[14][31] ) );
  DFFR_X1 \REGISTERS_reg[14][30]  ( .D(DATA_IN[30]), .CK(net18925), .RN(RST), 
        .Q(\REGISTERS[14][30] ) );
  DFFR_X1 \REGISTERS_reg[14][29]  ( .D(DATA_IN[29]), .CK(net18925), .RN(RST), 
        .Q(\REGISTERS[14][29] ) );
  DFFR_X1 \REGISTERS_reg[14][28]  ( .D(DATA_IN[28]), .CK(net18925), .RN(RST), 
        .Q(\REGISTERS[14][28] ) );
  DFFR_X1 \REGISTERS_reg[14][27]  ( .D(DATA_IN[27]), .CK(net18925), .RN(RST), 
        .Q(\REGISTERS[14][27] ) );
  DFFR_X1 \REGISTERS_reg[14][26]  ( .D(DATA_IN[26]), .CK(net18925), .RN(RST), 
        .Q(\REGISTERS[14][26] ) );
  DFFR_X1 \REGISTERS_reg[14][25]  ( .D(DATA_IN[25]), .CK(net18925), .RN(RST), 
        .Q(\REGISTERS[14][25] ) );
  DFFR_X1 \REGISTERS_reg[14][24]  ( .D(DATA_IN[24]), .CK(net18925), .RN(RST), 
        .Q(\REGISTERS[14][24] ) );
  DFFR_X1 \REGISTERS_reg[14][23]  ( .D(DATA_IN[23]), .CK(net18925), .RN(RST), 
        .Q(\REGISTERS[14][23] ) );
  DFFR_X1 \REGISTERS_reg[14][22]  ( .D(DATA_IN[22]), .CK(net18925), .RN(RST), 
        .Q(\REGISTERS[14][22] ) );
  DFFR_X1 \REGISTERS_reg[14][21]  ( .D(DATA_IN[21]), .CK(net18925), .RN(RST), 
        .Q(\REGISTERS[14][21] ) );
  DFFR_X1 \REGISTERS_reg[14][20]  ( .D(DATA_IN[20]), .CK(net18925), .RN(RST), 
        .Q(\REGISTERS[14][20] ) );
  DFFR_X1 \REGISTERS_reg[14][19]  ( .D(DATA_IN[19]), .CK(net18925), .RN(RST), 
        .Q(\REGISTERS[14][19] ) );
  DFFR_X1 \REGISTERS_reg[14][18]  ( .D(DATA_IN[18]), .CK(net18925), .RN(RST), 
        .Q(\REGISTERS[14][18] ) );
  DFFR_X1 \REGISTERS_reg[14][17]  ( .D(DATA_IN[17]), .CK(net18925), .RN(RST), 
        .Q(\REGISTERS[14][17] ) );
  DFFR_X1 \REGISTERS_reg[14][16]  ( .D(DATA_IN[16]), .CK(net18925), .RN(RST), 
        .Q(\REGISTERS[14][16] ) );
  DFFR_X1 \REGISTERS_reg[14][15]  ( .D(DATA_IN[15]), .CK(net18925), .RN(RST), 
        .Q(\REGISTERS[14][15] ) );
  DFFR_X1 \REGISTERS_reg[14][14]  ( .D(DATA_IN[14]), .CK(net18925), .RN(RST), 
        .Q(\REGISTERS[14][14] ) );
  DFFR_X1 \REGISTERS_reg[14][13]  ( .D(DATA_IN[13]), .CK(net18925), .RN(RST), 
        .Q(\REGISTERS[14][13] ) );
  DFFR_X1 \REGISTERS_reg[14][12]  ( .D(DATA_IN[12]), .CK(net18925), .RN(RST), 
        .Q(\REGISTERS[14][12] ) );
  DFFR_X1 \REGISTERS_reg[14][11]  ( .D(DATA_IN[11]), .CK(net18925), .RN(RST), 
        .Q(\REGISTERS[14][11] ) );
  DFFR_X1 \REGISTERS_reg[14][10]  ( .D(DATA_IN[10]), .CK(net18925), .RN(RST), 
        .Q(\REGISTERS[14][10] ) );
  DFFR_X1 \REGISTERS_reg[14][9]  ( .D(DATA_IN[9]), .CK(net18925), .RN(RST), 
        .Q(\REGISTERS[14][9] ) );
  DFFR_X1 \REGISTERS_reg[14][8]  ( .D(DATA_IN[8]), .CK(net18925), .RN(RST), 
        .Q(\REGISTERS[14][8] ) );
  DFFR_X1 \REGISTERS_reg[14][7]  ( .D(DATA_IN[7]), .CK(net18925), .RN(RST), 
        .Q(\REGISTERS[14][7] ) );
  DFFR_X1 \REGISTERS_reg[14][6]  ( .D(DATA_IN[6]), .CK(net18925), .RN(RST), 
        .Q(\REGISTERS[14][6] ) );
  DFFR_X1 \REGISTERS_reg[14][5]  ( .D(DATA_IN[5]), .CK(net18925), .RN(RST), 
        .Q(\REGISTERS[14][5] ) );
  DFFR_X1 \REGISTERS_reg[14][4]  ( .D(DATA_IN[4]), .CK(net18925), .RN(RST), 
        .Q(\REGISTERS[14][4] ) );
  DFFR_X1 \REGISTERS_reg[14][3]  ( .D(DATA_IN[3]), .CK(net18925), .RN(RST), 
        .Q(\REGISTERS[14][3] ) );
  DFFR_X1 \REGISTERS_reg[14][2]  ( .D(DATA_IN[2]), .CK(net18925), .RN(RST), 
        .Q(\REGISTERS[14][2] ) );
  DFFR_X1 \REGISTERS_reg[14][1]  ( .D(DATA_IN[1]), .CK(net18925), .RN(RST), 
        .Q(\REGISTERS[14][1] ) );
  DFFR_X1 \REGISTERS_reg[14][0]  ( .D(DATA_IN[0]), .CK(net18925), .RN(RST), 
        .Q(\REGISTERS[14][0] ) );
  DFFR_X1 \REGISTERS_reg[15][31]  ( .D(DATA_IN[31]), .CK(net18930), .RN(RST), 
        .Q(\REGISTERS[15][31] ) );
  DFFR_X1 \REGISTERS_reg[15][30]  ( .D(DATA_IN[30]), .CK(net18930), .RN(RST), 
        .Q(\REGISTERS[15][30] ) );
  DFFR_X1 \REGISTERS_reg[15][29]  ( .D(DATA_IN[29]), .CK(net18930), .RN(RST), 
        .Q(\REGISTERS[15][29] ) );
  DFFR_X1 \REGISTERS_reg[15][28]  ( .D(DATA_IN[28]), .CK(net18930), .RN(RST), 
        .Q(\REGISTERS[15][28] ) );
  DFFR_X1 \REGISTERS_reg[15][27]  ( .D(DATA_IN[27]), .CK(net18930), .RN(RST), 
        .Q(\REGISTERS[15][27] ) );
  DFFR_X1 \REGISTERS_reg[15][26]  ( .D(DATA_IN[26]), .CK(net18930), .RN(RST), 
        .Q(\REGISTERS[15][26] ) );
  DFFR_X1 \REGISTERS_reg[15][25]  ( .D(DATA_IN[25]), .CK(net18930), .RN(RST), 
        .Q(\REGISTERS[15][25] ) );
  DFFR_X1 \REGISTERS_reg[15][24]  ( .D(DATA_IN[24]), .CK(net18930), .RN(RST), 
        .Q(\REGISTERS[15][24] ) );
  DFFR_X1 \REGISTERS_reg[15][23]  ( .D(DATA_IN[23]), .CK(net18930), .RN(RST), 
        .Q(\REGISTERS[15][23] ) );
  DFFR_X1 \REGISTERS_reg[15][22]  ( .D(DATA_IN[22]), .CK(net18930), .RN(RST), 
        .Q(\REGISTERS[15][22] ) );
  DFFR_X1 \REGISTERS_reg[15][21]  ( .D(DATA_IN[21]), .CK(net18930), .RN(RST), 
        .Q(\REGISTERS[15][21] ) );
  DFFR_X1 \REGISTERS_reg[15][20]  ( .D(DATA_IN[20]), .CK(net18930), .RN(RST), 
        .Q(\REGISTERS[15][20] ) );
  DFFR_X1 \REGISTERS_reg[15][19]  ( .D(DATA_IN[19]), .CK(net18930), .RN(RST), 
        .Q(\REGISTERS[15][19] ) );
  DFFR_X1 \REGISTERS_reg[15][18]  ( .D(DATA_IN[18]), .CK(net18930), .RN(RST), 
        .Q(\REGISTERS[15][18] ) );
  DFFR_X1 \REGISTERS_reg[15][17]  ( .D(DATA_IN[17]), .CK(net18930), .RN(RST), 
        .Q(\REGISTERS[15][17] ) );
  DFFR_X1 \REGISTERS_reg[15][16]  ( .D(DATA_IN[16]), .CK(net18930), .RN(RST), 
        .Q(\REGISTERS[15][16] ) );
  DFFR_X1 \REGISTERS_reg[15][15]  ( .D(DATA_IN[15]), .CK(net18930), .RN(RST), 
        .Q(\REGISTERS[15][15] ) );
  DFFR_X1 \REGISTERS_reg[15][14]  ( .D(DATA_IN[14]), .CK(net18930), .RN(RST), 
        .Q(\REGISTERS[15][14] ) );
  DFFR_X1 \REGISTERS_reg[15][13]  ( .D(DATA_IN[13]), .CK(net18930), .RN(RST), 
        .Q(\REGISTERS[15][13] ) );
  DFFR_X1 \REGISTERS_reg[15][12]  ( .D(DATA_IN[12]), .CK(net18930), .RN(RST), 
        .Q(\REGISTERS[15][12] ) );
  DFFR_X1 \REGISTERS_reg[15][11]  ( .D(DATA_IN[11]), .CK(net18930), .RN(RST), 
        .Q(\REGISTERS[15][11] ) );
  DFFR_X1 \REGISTERS_reg[15][10]  ( .D(DATA_IN[10]), .CK(net18930), .RN(RST), 
        .Q(\REGISTERS[15][10] ) );
  DFFR_X1 \REGISTERS_reg[15][9]  ( .D(DATA_IN[9]), .CK(net18930), .RN(RST), 
        .Q(\REGISTERS[15][9] ) );
  DFFR_X1 \REGISTERS_reg[15][8]  ( .D(DATA_IN[8]), .CK(net18930), .RN(RST), 
        .Q(\REGISTERS[15][8] ) );
  DFFR_X1 \REGISTERS_reg[15][7]  ( .D(DATA_IN[7]), .CK(net18930), .RN(RST), 
        .Q(\REGISTERS[15][7] ) );
  DFFR_X1 \REGISTERS_reg[15][6]  ( .D(DATA_IN[6]), .CK(net18930), .RN(RST), 
        .Q(\REGISTERS[15][6] ) );
  DFFR_X1 \REGISTERS_reg[15][5]  ( .D(DATA_IN[5]), .CK(net18930), .RN(RST), 
        .Q(\REGISTERS[15][5] ) );
  DFFR_X1 \REGISTERS_reg[15][4]  ( .D(DATA_IN[4]), .CK(net18930), .RN(RST), 
        .Q(\REGISTERS[15][4] ) );
  DFFR_X1 \REGISTERS_reg[15][3]  ( .D(DATA_IN[3]), .CK(net18930), .RN(RST), 
        .Q(\REGISTERS[15][3] ) );
  DFFR_X1 \REGISTERS_reg[15][2]  ( .D(DATA_IN[2]), .CK(net18930), .RN(RST), 
        .Q(\REGISTERS[15][2] ) );
  DFFR_X1 \REGISTERS_reg[15][1]  ( .D(DATA_IN[1]), .CK(net18930), .RN(RST), 
        .Q(\REGISTERS[15][1] ) );
  DFFR_X1 \REGISTERS_reg[15][0]  ( .D(DATA_IN[0]), .CK(net18930), .RN(RST), 
        .Q(\REGISTERS[15][0] ) );
  DFFR_X1 \REGISTERS_reg[16][31]  ( .D(DATA_IN[31]), .CK(net18935), .RN(RST), 
        .Q(\REGISTERS[16][31] ) );
  DFFR_X1 \REGISTERS_reg[16][30]  ( .D(DATA_IN[30]), .CK(net18935), .RN(RST), 
        .Q(\REGISTERS[16][30] ) );
  DFFR_X1 \REGISTERS_reg[16][29]  ( .D(DATA_IN[29]), .CK(net18935), .RN(RST), 
        .Q(\REGISTERS[16][29] ) );
  DFFR_X1 \REGISTERS_reg[16][28]  ( .D(DATA_IN[28]), .CK(net18935), .RN(RST), 
        .Q(\REGISTERS[16][28] ) );
  DFFR_X1 \REGISTERS_reg[16][27]  ( .D(DATA_IN[27]), .CK(net18935), .RN(RST), 
        .Q(\REGISTERS[16][27] ) );
  DFFR_X1 \REGISTERS_reg[16][26]  ( .D(DATA_IN[26]), .CK(net18935), .RN(RST), 
        .Q(\REGISTERS[16][26] ) );
  DFFR_X1 \REGISTERS_reg[16][25]  ( .D(DATA_IN[25]), .CK(net18935), .RN(RST), 
        .Q(\REGISTERS[16][25] ) );
  DFFR_X1 \REGISTERS_reg[16][24]  ( .D(DATA_IN[24]), .CK(net18935), .RN(RST), 
        .Q(\REGISTERS[16][24] ) );
  DFFR_X1 \REGISTERS_reg[16][23]  ( .D(DATA_IN[23]), .CK(net18935), .RN(RST), 
        .Q(\REGISTERS[16][23] ) );
  DFFR_X1 \REGISTERS_reg[16][22]  ( .D(DATA_IN[22]), .CK(net18935), .RN(RST), 
        .Q(\REGISTERS[16][22] ) );
  DFFR_X1 \REGISTERS_reg[16][21]  ( .D(DATA_IN[21]), .CK(net18935), .RN(RST), 
        .Q(\REGISTERS[16][21] ) );
  DFFR_X1 \REGISTERS_reg[16][20]  ( .D(DATA_IN[20]), .CK(net18935), .RN(RST), 
        .Q(\REGISTERS[16][20] ) );
  DFFR_X1 \REGISTERS_reg[16][19]  ( .D(DATA_IN[19]), .CK(net18935), .RN(RST), 
        .Q(\REGISTERS[16][19] ) );
  DFFR_X1 \REGISTERS_reg[16][18]  ( .D(DATA_IN[18]), .CK(net18935), .RN(RST), 
        .Q(\REGISTERS[16][18] ) );
  DFFR_X1 \REGISTERS_reg[16][17]  ( .D(DATA_IN[17]), .CK(net18935), .RN(RST), 
        .Q(\REGISTERS[16][17] ) );
  DFFR_X1 \REGISTERS_reg[16][16]  ( .D(DATA_IN[16]), .CK(net18935), .RN(RST), 
        .Q(\REGISTERS[16][16] ) );
  DFFR_X1 \REGISTERS_reg[16][15]  ( .D(DATA_IN[15]), .CK(net18935), .RN(RST), 
        .Q(\REGISTERS[16][15] ) );
  DFFR_X1 \REGISTERS_reg[16][14]  ( .D(DATA_IN[14]), .CK(net18935), .RN(RST), 
        .Q(\REGISTERS[16][14] ) );
  DFFR_X1 \REGISTERS_reg[16][13]  ( .D(DATA_IN[13]), .CK(net18935), .RN(RST), 
        .Q(\REGISTERS[16][13] ) );
  DFFR_X1 \REGISTERS_reg[16][12]  ( .D(DATA_IN[12]), .CK(net18935), .RN(RST), 
        .Q(\REGISTERS[16][12] ) );
  DFFR_X1 \REGISTERS_reg[16][11]  ( .D(DATA_IN[11]), .CK(net18935), .RN(RST), 
        .Q(\REGISTERS[16][11] ) );
  DFFR_X1 \REGISTERS_reg[16][10]  ( .D(DATA_IN[10]), .CK(net18935), .RN(RST), 
        .Q(\REGISTERS[16][10] ) );
  DFFR_X1 \REGISTERS_reg[16][9]  ( .D(DATA_IN[9]), .CK(net18935), .RN(RST), 
        .Q(\REGISTERS[16][9] ) );
  DFFR_X1 \REGISTERS_reg[16][8]  ( .D(DATA_IN[8]), .CK(net18935), .RN(RST), 
        .Q(\REGISTERS[16][8] ) );
  DFFR_X1 \REGISTERS_reg[16][7]  ( .D(DATA_IN[7]), .CK(net18935), .RN(RST), 
        .Q(\REGISTERS[16][7] ) );
  DFFR_X1 \REGISTERS_reg[16][6]  ( .D(DATA_IN[6]), .CK(net18935), .RN(RST), 
        .Q(\REGISTERS[16][6] ) );
  DFFR_X1 \REGISTERS_reg[16][5]  ( .D(DATA_IN[5]), .CK(net18935), .RN(RST), 
        .Q(\REGISTERS[16][5] ) );
  DFFR_X1 \REGISTERS_reg[16][4]  ( .D(DATA_IN[4]), .CK(net18935), .RN(RST), 
        .Q(\REGISTERS[16][4] ) );
  DFFR_X1 \REGISTERS_reg[16][3]  ( .D(DATA_IN[3]), .CK(net18935), .RN(RST), 
        .Q(\REGISTERS[16][3] ) );
  DFFR_X1 \REGISTERS_reg[16][2]  ( .D(DATA_IN[2]), .CK(net18935), .RN(RST), 
        .Q(\REGISTERS[16][2] ) );
  DFFR_X1 \REGISTERS_reg[16][1]  ( .D(DATA_IN[1]), .CK(net18935), .RN(RST), 
        .Q(\REGISTERS[16][1] ) );
  DFFR_X1 \REGISTERS_reg[16][0]  ( .D(DATA_IN[0]), .CK(net18935), .RN(RST), 
        .Q(\REGISTERS[16][0] ) );
  DFFR_X1 \REGISTERS_reg[17][31]  ( .D(DATA_IN[31]), .CK(net18940), .RN(RST), 
        .Q(\REGISTERS[17][31] ) );
  DFFR_X1 \REGISTERS_reg[17][30]  ( .D(DATA_IN[30]), .CK(net18940), .RN(RST), 
        .Q(\REGISTERS[17][30] ) );
  DFFR_X1 \REGISTERS_reg[17][29]  ( .D(DATA_IN[29]), .CK(net18940), .RN(RST), 
        .Q(\REGISTERS[17][29] ) );
  DFFR_X1 \REGISTERS_reg[17][28]  ( .D(DATA_IN[28]), .CK(net18940), .RN(RST), 
        .Q(\REGISTERS[17][28] ) );
  DFFR_X1 \REGISTERS_reg[17][27]  ( .D(DATA_IN[27]), .CK(net18940), .RN(RST), 
        .Q(\REGISTERS[17][27] ) );
  DFFR_X1 \REGISTERS_reg[17][26]  ( .D(DATA_IN[26]), .CK(net18940), .RN(RST), 
        .Q(\REGISTERS[17][26] ) );
  DFFR_X1 \REGISTERS_reg[17][25]  ( .D(DATA_IN[25]), .CK(net18940), .RN(RST), 
        .Q(\REGISTERS[17][25] ) );
  DFFR_X1 \REGISTERS_reg[17][24]  ( .D(DATA_IN[24]), .CK(net18940), .RN(RST), 
        .Q(\REGISTERS[17][24] ) );
  DFFR_X1 \REGISTERS_reg[17][23]  ( .D(DATA_IN[23]), .CK(net18940), .RN(RST), 
        .Q(\REGISTERS[17][23] ) );
  DFFR_X1 \REGISTERS_reg[17][22]  ( .D(DATA_IN[22]), .CK(net18940), .RN(RST), 
        .Q(\REGISTERS[17][22] ) );
  DFFR_X1 \REGISTERS_reg[17][21]  ( .D(DATA_IN[21]), .CK(net18940), .RN(RST), 
        .Q(\REGISTERS[17][21] ) );
  DFFR_X1 \REGISTERS_reg[17][20]  ( .D(DATA_IN[20]), .CK(net18940), .RN(RST), 
        .Q(\REGISTERS[17][20] ) );
  DFFR_X1 \REGISTERS_reg[17][19]  ( .D(DATA_IN[19]), .CK(net18940), .RN(RST), 
        .Q(\REGISTERS[17][19] ) );
  DFFR_X1 \REGISTERS_reg[17][18]  ( .D(DATA_IN[18]), .CK(net18940), .RN(RST), 
        .Q(\REGISTERS[17][18] ) );
  DFFR_X1 \REGISTERS_reg[17][17]  ( .D(DATA_IN[17]), .CK(net18940), .RN(RST), 
        .Q(\REGISTERS[17][17] ) );
  DFFR_X1 \REGISTERS_reg[17][16]  ( .D(DATA_IN[16]), .CK(net18940), .RN(RST), 
        .Q(\REGISTERS[17][16] ) );
  DFFR_X1 \REGISTERS_reg[17][15]  ( .D(DATA_IN[15]), .CK(net18940), .RN(RST), 
        .Q(\REGISTERS[17][15] ) );
  DFFR_X1 \REGISTERS_reg[17][14]  ( .D(DATA_IN[14]), .CK(net18940), .RN(RST), 
        .Q(\REGISTERS[17][14] ) );
  DFFR_X1 \REGISTERS_reg[17][13]  ( .D(DATA_IN[13]), .CK(net18940), .RN(RST), 
        .Q(\REGISTERS[17][13] ) );
  DFFR_X1 \REGISTERS_reg[17][12]  ( .D(DATA_IN[12]), .CK(net18940), .RN(RST), 
        .Q(\REGISTERS[17][12] ) );
  DFFR_X1 \REGISTERS_reg[17][11]  ( .D(DATA_IN[11]), .CK(net18940), .RN(RST), 
        .Q(\REGISTERS[17][11] ) );
  DFFR_X1 \REGISTERS_reg[17][10]  ( .D(DATA_IN[10]), .CK(net18940), .RN(RST), 
        .Q(\REGISTERS[17][10] ) );
  DFFR_X1 \REGISTERS_reg[17][9]  ( .D(DATA_IN[9]), .CK(net18940), .RN(RST), 
        .Q(\REGISTERS[17][9] ) );
  DFFR_X1 \REGISTERS_reg[17][8]  ( .D(DATA_IN[8]), .CK(net18940), .RN(RST), 
        .Q(\REGISTERS[17][8] ) );
  DFFR_X1 \REGISTERS_reg[17][7]  ( .D(DATA_IN[7]), .CK(net18940), .RN(RST), 
        .Q(\REGISTERS[17][7] ) );
  DFFR_X1 \REGISTERS_reg[17][6]  ( .D(DATA_IN[6]), .CK(net18940), .RN(RST), 
        .Q(\REGISTERS[17][6] ) );
  DFFR_X1 \REGISTERS_reg[17][5]  ( .D(DATA_IN[5]), .CK(net18940), .RN(RST), 
        .Q(\REGISTERS[17][5] ) );
  DFFR_X1 \REGISTERS_reg[17][4]  ( .D(DATA_IN[4]), .CK(net18940), .RN(RST), 
        .Q(\REGISTERS[17][4] ) );
  DFFR_X1 \REGISTERS_reg[17][3]  ( .D(DATA_IN[3]), .CK(net18940), .RN(RST), 
        .Q(\REGISTERS[17][3] ) );
  DFFR_X1 \REGISTERS_reg[17][2]  ( .D(DATA_IN[2]), .CK(net18940), .RN(RST), 
        .Q(\REGISTERS[17][2] ) );
  DFFR_X1 \REGISTERS_reg[17][1]  ( .D(DATA_IN[1]), .CK(net18940), .RN(RST), 
        .Q(\REGISTERS[17][1] ) );
  DFFR_X1 \REGISTERS_reg[17][0]  ( .D(DATA_IN[0]), .CK(net18940), .RN(RST), 
        .Q(\REGISTERS[17][0] ) );
  DFFR_X1 \REGISTERS_reg[18][31]  ( .D(DATA_IN[31]), .CK(net18945), .RN(RST), 
        .Q(\REGISTERS[18][31] ) );
  DFFR_X1 \REGISTERS_reg[18][30]  ( .D(DATA_IN[30]), .CK(net18945), .RN(RST), 
        .Q(\REGISTERS[18][30] ) );
  DFFR_X1 \REGISTERS_reg[18][29]  ( .D(DATA_IN[29]), .CK(net18945), .RN(RST), 
        .Q(\REGISTERS[18][29] ) );
  DFFR_X1 \REGISTERS_reg[18][28]  ( .D(DATA_IN[28]), .CK(net18945), .RN(RST), 
        .Q(\REGISTERS[18][28] ) );
  DFFR_X1 \REGISTERS_reg[18][27]  ( .D(DATA_IN[27]), .CK(net18945), .RN(RST), 
        .Q(\REGISTERS[18][27] ) );
  DFFR_X1 \REGISTERS_reg[18][26]  ( .D(DATA_IN[26]), .CK(net18945), .RN(RST), 
        .Q(\REGISTERS[18][26] ) );
  DFFR_X1 \REGISTERS_reg[18][25]  ( .D(DATA_IN[25]), .CK(net18945), .RN(RST), 
        .Q(\REGISTERS[18][25] ) );
  DFFR_X1 \REGISTERS_reg[18][24]  ( .D(DATA_IN[24]), .CK(net18945), .RN(RST), 
        .Q(\REGISTERS[18][24] ) );
  DFFR_X1 \REGISTERS_reg[18][23]  ( .D(DATA_IN[23]), .CK(net18945), .RN(RST), 
        .Q(\REGISTERS[18][23] ) );
  DFFR_X1 \REGISTERS_reg[18][22]  ( .D(DATA_IN[22]), .CK(net18945), .RN(RST), 
        .Q(\REGISTERS[18][22] ) );
  DFFR_X1 \REGISTERS_reg[18][21]  ( .D(DATA_IN[21]), .CK(net18945), .RN(RST), 
        .Q(\REGISTERS[18][21] ) );
  DFFR_X1 \REGISTERS_reg[18][20]  ( .D(DATA_IN[20]), .CK(net18945), .RN(RST), 
        .Q(\REGISTERS[18][20] ) );
  DFFR_X1 \REGISTERS_reg[18][19]  ( .D(DATA_IN[19]), .CK(net18945), .RN(RST), 
        .Q(\REGISTERS[18][19] ) );
  DFFR_X1 \REGISTERS_reg[18][18]  ( .D(DATA_IN[18]), .CK(net18945), .RN(RST), 
        .Q(\REGISTERS[18][18] ) );
  DFFR_X1 \REGISTERS_reg[18][17]  ( .D(DATA_IN[17]), .CK(net18945), .RN(RST), 
        .Q(\REGISTERS[18][17] ) );
  DFFR_X1 \REGISTERS_reg[18][16]  ( .D(DATA_IN[16]), .CK(net18945), .RN(RST), 
        .Q(\REGISTERS[18][16] ) );
  DFFR_X1 \REGISTERS_reg[18][15]  ( .D(DATA_IN[15]), .CK(net18945), .RN(RST), 
        .Q(\REGISTERS[18][15] ) );
  DFFR_X1 \REGISTERS_reg[18][14]  ( .D(DATA_IN[14]), .CK(net18945), .RN(RST), 
        .Q(\REGISTERS[18][14] ) );
  DFFR_X1 \REGISTERS_reg[18][13]  ( .D(DATA_IN[13]), .CK(net18945), .RN(RST), 
        .Q(\REGISTERS[18][13] ) );
  DFFR_X1 \REGISTERS_reg[18][12]  ( .D(DATA_IN[12]), .CK(net18945), .RN(RST), 
        .Q(\REGISTERS[18][12] ) );
  DFFR_X1 \REGISTERS_reg[18][11]  ( .D(DATA_IN[11]), .CK(net18945), .RN(RST), 
        .Q(\REGISTERS[18][11] ) );
  DFFR_X1 \REGISTERS_reg[18][10]  ( .D(DATA_IN[10]), .CK(net18945), .RN(RST), 
        .Q(\REGISTERS[18][10] ) );
  DFFR_X1 \REGISTERS_reg[18][9]  ( .D(DATA_IN[9]), .CK(net18945), .RN(RST), 
        .Q(\REGISTERS[18][9] ) );
  DFFR_X1 \REGISTERS_reg[18][8]  ( .D(DATA_IN[8]), .CK(net18945), .RN(RST), 
        .Q(\REGISTERS[18][8] ) );
  DFFR_X1 \REGISTERS_reg[18][7]  ( .D(DATA_IN[7]), .CK(net18945), .RN(RST), 
        .Q(\REGISTERS[18][7] ) );
  DFFR_X1 \REGISTERS_reg[18][6]  ( .D(DATA_IN[6]), .CK(net18945), .RN(RST), 
        .Q(\REGISTERS[18][6] ) );
  DFFR_X1 \REGISTERS_reg[18][5]  ( .D(DATA_IN[5]), .CK(net18945), .RN(RST), 
        .Q(\REGISTERS[18][5] ) );
  DFFR_X1 \REGISTERS_reg[18][4]  ( .D(DATA_IN[4]), .CK(net18945), .RN(RST), 
        .Q(\REGISTERS[18][4] ) );
  DFFR_X1 \REGISTERS_reg[18][3]  ( .D(DATA_IN[3]), .CK(net18945), .RN(RST), 
        .Q(\REGISTERS[18][3] ) );
  DFFR_X1 \REGISTERS_reg[18][2]  ( .D(DATA_IN[2]), .CK(net18945), .RN(RST), 
        .Q(\REGISTERS[18][2] ) );
  DFFR_X1 \REGISTERS_reg[18][1]  ( .D(DATA_IN[1]), .CK(net18945), .RN(RST), 
        .Q(\REGISTERS[18][1] ) );
  DFFR_X1 \REGISTERS_reg[18][0]  ( .D(DATA_IN[0]), .CK(net18945), .RN(RST), 
        .Q(\REGISTERS[18][0] ) );
  DFFR_X1 \REGISTERS_reg[19][31]  ( .D(DATA_IN[31]), .CK(net18950), .RN(RST), 
        .Q(\REGISTERS[19][31] ) );
  DFFR_X1 \REGISTERS_reg[19][30]  ( .D(DATA_IN[30]), .CK(net18950), .RN(RST), 
        .Q(\REGISTERS[19][30] ) );
  DFFR_X1 \REGISTERS_reg[19][29]  ( .D(DATA_IN[29]), .CK(net18950), .RN(RST), 
        .Q(\REGISTERS[19][29] ) );
  DFFR_X1 \REGISTERS_reg[19][28]  ( .D(DATA_IN[28]), .CK(net18950), .RN(RST), 
        .Q(\REGISTERS[19][28] ) );
  DFFR_X1 \REGISTERS_reg[19][27]  ( .D(DATA_IN[27]), .CK(net18950), .RN(RST), 
        .Q(\REGISTERS[19][27] ) );
  DFFR_X1 \REGISTERS_reg[19][26]  ( .D(DATA_IN[26]), .CK(net18950), .RN(RST), 
        .Q(\REGISTERS[19][26] ) );
  DFFR_X1 \REGISTERS_reg[19][25]  ( .D(DATA_IN[25]), .CK(net18950), .RN(RST), 
        .Q(\REGISTERS[19][25] ) );
  DFFR_X1 \REGISTERS_reg[19][24]  ( .D(DATA_IN[24]), .CK(net18950), .RN(RST), 
        .Q(\REGISTERS[19][24] ) );
  DFFR_X1 \REGISTERS_reg[19][23]  ( .D(DATA_IN[23]), .CK(net18950), .RN(RST), 
        .Q(\REGISTERS[19][23] ) );
  DFFR_X1 \REGISTERS_reg[19][22]  ( .D(DATA_IN[22]), .CK(net18950), .RN(RST), 
        .Q(\REGISTERS[19][22] ) );
  DFFR_X1 \REGISTERS_reg[19][21]  ( .D(DATA_IN[21]), .CK(net18950), .RN(RST), 
        .Q(\REGISTERS[19][21] ) );
  DFFR_X1 \REGISTERS_reg[19][20]  ( .D(DATA_IN[20]), .CK(net18950), .RN(RST), 
        .Q(\REGISTERS[19][20] ) );
  DFFR_X1 \REGISTERS_reg[19][19]  ( .D(DATA_IN[19]), .CK(net18950), .RN(RST), 
        .Q(\REGISTERS[19][19] ) );
  DFFR_X1 \REGISTERS_reg[19][18]  ( .D(DATA_IN[18]), .CK(net18950), .RN(RST), 
        .Q(\REGISTERS[19][18] ) );
  DFFR_X1 \REGISTERS_reg[19][17]  ( .D(DATA_IN[17]), .CK(net18950), .RN(RST), 
        .Q(\REGISTERS[19][17] ) );
  DFFR_X1 \REGISTERS_reg[19][16]  ( .D(DATA_IN[16]), .CK(net18950), .RN(RST), 
        .Q(\REGISTERS[19][16] ) );
  DFFR_X1 \REGISTERS_reg[19][15]  ( .D(DATA_IN[15]), .CK(net18950), .RN(RST), 
        .Q(\REGISTERS[19][15] ) );
  DFFR_X1 \REGISTERS_reg[19][14]  ( .D(DATA_IN[14]), .CK(net18950), .RN(RST), 
        .Q(\REGISTERS[19][14] ) );
  DFFR_X1 \REGISTERS_reg[19][13]  ( .D(DATA_IN[13]), .CK(net18950), .RN(RST), 
        .Q(\REGISTERS[19][13] ) );
  DFFR_X1 \REGISTERS_reg[19][12]  ( .D(DATA_IN[12]), .CK(net18950), .RN(RST), 
        .Q(\REGISTERS[19][12] ) );
  DFFR_X1 \REGISTERS_reg[19][11]  ( .D(DATA_IN[11]), .CK(net18950), .RN(RST), 
        .Q(\REGISTERS[19][11] ) );
  DFFR_X1 \REGISTERS_reg[19][10]  ( .D(DATA_IN[10]), .CK(net18950), .RN(RST), 
        .Q(\REGISTERS[19][10] ) );
  DFFR_X1 \REGISTERS_reg[19][9]  ( .D(DATA_IN[9]), .CK(net18950), .RN(RST), 
        .Q(\REGISTERS[19][9] ) );
  DFFR_X1 \REGISTERS_reg[19][8]  ( .D(DATA_IN[8]), .CK(net18950), .RN(RST), 
        .Q(\REGISTERS[19][8] ) );
  DFFR_X1 \REGISTERS_reg[19][7]  ( .D(DATA_IN[7]), .CK(net18950), .RN(RST), 
        .Q(\REGISTERS[19][7] ) );
  DFFR_X1 \REGISTERS_reg[19][6]  ( .D(DATA_IN[6]), .CK(net18950), .RN(RST), 
        .Q(\REGISTERS[19][6] ) );
  DFFR_X1 \REGISTERS_reg[19][5]  ( .D(DATA_IN[5]), .CK(net18950), .RN(RST), 
        .Q(\REGISTERS[19][5] ) );
  DFFR_X1 \REGISTERS_reg[19][4]  ( .D(DATA_IN[4]), .CK(net18950), .RN(RST), 
        .Q(\REGISTERS[19][4] ) );
  DFFR_X1 \REGISTERS_reg[19][3]  ( .D(DATA_IN[3]), .CK(net18950), .RN(RST), 
        .Q(\REGISTERS[19][3] ) );
  DFFR_X1 \REGISTERS_reg[19][2]  ( .D(DATA_IN[2]), .CK(net18950), .RN(RST), 
        .Q(\REGISTERS[19][2] ) );
  DFFR_X1 \REGISTERS_reg[19][1]  ( .D(DATA_IN[1]), .CK(net18950), .RN(RST), 
        .Q(\REGISTERS[19][1] ) );
  DFFR_X1 \REGISTERS_reg[19][0]  ( .D(DATA_IN[0]), .CK(net18950), .RN(RST), 
        .Q(\REGISTERS[19][0] ) );
  DFFR_X1 \REGISTERS_reg[20][31]  ( .D(DATA_IN[31]), .CK(net18955), .RN(RST), 
        .Q(\REGISTERS[20][31] ) );
  DFFR_X1 \REGISTERS_reg[20][30]  ( .D(DATA_IN[30]), .CK(net18955), .RN(RST), 
        .Q(\REGISTERS[20][30] ) );
  DFFR_X1 \REGISTERS_reg[20][29]  ( .D(DATA_IN[29]), .CK(net18955), .RN(RST), 
        .Q(\REGISTERS[20][29] ) );
  DFFR_X1 \REGISTERS_reg[20][28]  ( .D(DATA_IN[28]), .CK(net18955), .RN(RST), 
        .Q(\REGISTERS[20][28] ) );
  DFFR_X1 \REGISTERS_reg[20][27]  ( .D(DATA_IN[27]), .CK(net18955), .RN(RST), 
        .Q(\REGISTERS[20][27] ) );
  DFFR_X1 \REGISTERS_reg[20][26]  ( .D(DATA_IN[26]), .CK(net18955), .RN(RST), 
        .Q(\REGISTERS[20][26] ) );
  DFFR_X1 \REGISTERS_reg[20][25]  ( .D(DATA_IN[25]), .CK(net18955), .RN(RST), 
        .Q(\REGISTERS[20][25] ) );
  DFFR_X1 \REGISTERS_reg[20][24]  ( .D(DATA_IN[24]), .CK(net18955), .RN(RST), 
        .Q(\REGISTERS[20][24] ) );
  DFFR_X1 \REGISTERS_reg[20][23]  ( .D(DATA_IN[23]), .CK(net18955), .RN(RST), 
        .Q(\REGISTERS[20][23] ) );
  DFFR_X1 \REGISTERS_reg[20][22]  ( .D(DATA_IN[22]), .CK(net18955), .RN(RST), 
        .Q(\REGISTERS[20][22] ) );
  DFFR_X1 \REGISTERS_reg[20][21]  ( .D(DATA_IN[21]), .CK(net18955), .RN(RST), 
        .Q(\REGISTERS[20][21] ) );
  DFFR_X1 \REGISTERS_reg[20][20]  ( .D(DATA_IN[20]), .CK(net18955), .RN(RST), 
        .Q(\REGISTERS[20][20] ) );
  DFFR_X1 \REGISTERS_reg[20][19]  ( .D(DATA_IN[19]), .CK(net18955), .RN(RST), 
        .Q(\REGISTERS[20][19] ) );
  DFFR_X1 \REGISTERS_reg[20][18]  ( .D(DATA_IN[18]), .CK(net18955), .RN(RST), 
        .Q(\REGISTERS[20][18] ) );
  DFFR_X1 \REGISTERS_reg[20][17]  ( .D(DATA_IN[17]), .CK(net18955), .RN(RST), 
        .Q(\REGISTERS[20][17] ) );
  DFFR_X1 \REGISTERS_reg[20][16]  ( .D(DATA_IN[16]), .CK(net18955), .RN(RST), 
        .Q(\REGISTERS[20][16] ) );
  DFFR_X1 \REGISTERS_reg[20][15]  ( .D(DATA_IN[15]), .CK(net18955), .RN(RST), 
        .Q(\REGISTERS[20][15] ) );
  DFFR_X1 \REGISTERS_reg[20][14]  ( .D(DATA_IN[14]), .CK(net18955), .RN(RST), 
        .Q(\REGISTERS[20][14] ) );
  DFFR_X1 \REGISTERS_reg[20][13]  ( .D(DATA_IN[13]), .CK(net18955), .RN(RST), 
        .Q(\REGISTERS[20][13] ) );
  DFFR_X1 \REGISTERS_reg[20][12]  ( .D(DATA_IN[12]), .CK(net18955), .RN(RST), 
        .Q(\REGISTERS[20][12] ) );
  DFFR_X1 \REGISTERS_reg[20][11]  ( .D(DATA_IN[11]), .CK(net18955), .RN(RST), 
        .Q(\REGISTERS[20][11] ) );
  DFFR_X1 \REGISTERS_reg[20][10]  ( .D(DATA_IN[10]), .CK(net18955), .RN(RST), 
        .Q(\REGISTERS[20][10] ) );
  DFFR_X1 \REGISTERS_reg[20][9]  ( .D(DATA_IN[9]), .CK(net18955), .RN(RST), 
        .Q(\REGISTERS[20][9] ) );
  DFFR_X1 \REGISTERS_reg[20][8]  ( .D(DATA_IN[8]), .CK(net18955), .RN(RST), 
        .Q(\REGISTERS[20][8] ) );
  DFFR_X1 \REGISTERS_reg[20][7]  ( .D(DATA_IN[7]), .CK(net18955), .RN(RST), 
        .Q(\REGISTERS[20][7] ) );
  DFFR_X1 \REGISTERS_reg[20][6]  ( .D(DATA_IN[6]), .CK(net18955), .RN(RST), 
        .Q(\REGISTERS[20][6] ) );
  DFFR_X1 \REGISTERS_reg[20][5]  ( .D(DATA_IN[5]), .CK(net18955), .RN(RST), 
        .Q(\REGISTERS[20][5] ) );
  DFFR_X1 \REGISTERS_reg[20][4]  ( .D(DATA_IN[4]), .CK(net18955), .RN(RST), 
        .Q(\REGISTERS[20][4] ) );
  DFFR_X1 \REGISTERS_reg[20][3]  ( .D(DATA_IN[3]), .CK(net18955), .RN(RST), 
        .Q(\REGISTERS[20][3] ) );
  DFFR_X1 \REGISTERS_reg[20][2]  ( .D(DATA_IN[2]), .CK(net18955), .RN(RST), 
        .Q(\REGISTERS[20][2] ) );
  DFFR_X1 \REGISTERS_reg[20][1]  ( .D(DATA_IN[1]), .CK(net18955), .RN(RST), 
        .Q(\REGISTERS[20][1] ) );
  DFFR_X1 \REGISTERS_reg[20][0]  ( .D(DATA_IN[0]), .CK(net18955), .RN(RST), 
        .Q(\REGISTERS[20][0] ) );
  DFFR_X1 \REGISTERS_reg[21][31]  ( .D(DATA_IN[31]), .CK(net18960), .RN(RST), 
        .Q(\REGISTERS[21][31] ) );
  DFFR_X1 \REGISTERS_reg[21][30]  ( .D(DATA_IN[30]), .CK(net18960), .RN(RST), 
        .Q(\REGISTERS[21][30] ) );
  DFFR_X1 \REGISTERS_reg[21][29]  ( .D(DATA_IN[29]), .CK(net18960), .RN(RST), 
        .Q(\REGISTERS[21][29] ) );
  DFFR_X1 \REGISTERS_reg[21][28]  ( .D(DATA_IN[28]), .CK(net18960), .RN(RST), 
        .Q(\REGISTERS[21][28] ) );
  DFFR_X1 \REGISTERS_reg[21][27]  ( .D(DATA_IN[27]), .CK(net18960), .RN(RST), 
        .Q(\REGISTERS[21][27] ) );
  DFFR_X1 \REGISTERS_reg[21][26]  ( .D(DATA_IN[26]), .CK(net18960), .RN(RST), 
        .Q(\REGISTERS[21][26] ) );
  DFFR_X1 \REGISTERS_reg[21][25]  ( .D(DATA_IN[25]), .CK(net18960), .RN(RST), 
        .Q(\REGISTERS[21][25] ) );
  DFFR_X1 \REGISTERS_reg[21][24]  ( .D(DATA_IN[24]), .CK(net18960), .RN(RST), 
        .Q(\REGISTERS[21][24] ) );
  DFFR_X1 \REGISTERS_reg[21][23]  ( .D(DATA_IN[23]), .CK(net18960), .RN(RST), 
        .Q(\REGISTERS[21][23] ) );
  DFFR_X1 \REGISTERS_reg[21][22]  ( .D(DATA_IN[22]), .CK(net18960), .RN(RST), 
        .Q(\REGISTERS[21][22] ) );
  DFFR_X1 \REGISTERS_reg[21][21]  ( .D(DATA_IN[21]), .CK(net18960), .RN(RST), 
        .Q(\REGISTERS[21][21] ) );
  DFFR_X1 \REGISTERS_reg[21][20]  ( .D(DATA_IN[20]), .CK(net18960), .RN(RST), 
        .Q(\REGISTERS[21][20] ) );
  DFFR_X1 \REGISTERS_reg[21][19]  ( .D(DATA_IN[19]), .CK(net18960), .RN(RST), 
        .Q(\REGISTERS[21][19] ) );
  DFFR_X1 \REGISTERS_reg[21][18]  ( .D(DATA_IN[18]), .CK(net18960), .RN(RST), 
        .Q(\REGISTERS[21][18] ) );
  DFFR_X1 \REGISTERS_reg[21][17]  ( .D(DATA_IN[17]), .CK(net18960), .RN(RST), 
        .Q(\REGISTERS[21][17] ) );
  DFFR_X1 \REGISTERS_reg[21][16]  ( .D(DATA_IN[16]), .CK(net18960), .RN(RST), 
        .Q(\REGISTERS[21][16] ) );
  DFFR_X1 \REGISTERS_reg[21][15]  ( .D(DATA_IN[15]), .CK(net18960), .RN(RST), 
        .Q(\REGISTERS[21][15] ) );
  DFFR_X1 \REGISTERS_reg[21][14]  ( .D(DATA_IN[14]), .CK(net18960), .RN(RST), 
        .Q(\REGISTERS[21][14] ) );
  DFFR_X1 \REGISTERS_reg[21][13]  ( .D(DATA_IN[13]), .CK(net18960), .RN(RST), 
        .Q(\REGISTERS[21][13] ) );
  DFFR_X1 \REGISTERS_reg[21][12]  ( .D(DATA_IN[12]), .CK(net18960), .RN(RST), 
        .Q(\REGISTERS[21][12] ) );
  DFFR_X1 \REGISTERS_reg[21][11]  ( .D(DATA_IN[11]), .CK(net18960), .RN(RST), 
        .Q(\REGISTERS[21][11] ) );
  DFFR_X1 \REGISTERS_reg[21][10]  ( .D(DATA_IN[10]), .CK(net18960), .RN(RST), 
        .Q(\REGISTERS[21][10] ) );
  DFFR_X1 \REGISTERS_reg[21][9]  ( .D(DATA_IN[9]), .CK(net18960), .RN(RST), 
        .Q(\REGISTERS[21][9] ) );
  DFFR_X1 \REGISTERS_reg[21][8]  ( .D(DATA_IN[8]), .CK(net18960), .RN(RST), 
        .Q(\REGISTERS[21][8] ) );
  DFFR_X1 \REGISTERS_reg[21][7]  ( .D(DATA_IN[7]), .CK(net18960), .RN(RST), 
        .Q(\REGISTERS[21][7] ) );
  DFFR_X1 \REGISTERS_reg[21][6]  ( .D(DATA_IN[6]), .CK(net18960), .RN(RST), 
        .Q(\REGISTERS[21][6] ) );
  DFFR_X1 \REGISTERS_reg[21][5]  ( .D(DATA_IN[5]), .CK(net18960), .RN(RST), 
        .Q(\REGISTERS[21][5] ) );
  DFFR_X1 \REGISTERS_reg[21][4]  ( .D(DATA_IN[4]), .CK(net18960), .RN(RST), 
        .Q(\REGISTERS[21][4] ) );
  DFFR_X1 \REGISTERS_reg[21][3]  ( .D(DATA_IN[3]), .CK(net18960), .RN(RST), 
        .Q(\REGISTERS[21][3] ) );
  DFFR_X1 \REGISTERS_reg[21][2]  ( .D(DATA_IN[2]), .CK(net18960), .RN(RST), 
        .Q(\REGISTERS[21][2] ) );
  DFFR_X1 \REGISTERS_reg[21][1]  ( .D(DATA_IN[1]), .CK(net18960), .RN(RST), 
        .Q(\REGISTERS[21][1] ) );
  DFFR_X1 \REGISTERS_reg[21][0]  ( .D(DATA_IN[0]), .CK(net18960), .RN(RST), 
        .Q(\REGISTERS[21][0] ) );
  DFFR_X1 \REGISTERS_reg[22][31]  ( .D(DATA_IN[31]), .CK(net18965), .RN(RST), 
        .Q(\REGISTERS[22][31] ) );
  DFFR_X1 \REGISTERS_reg[22][30]  ( .D(DATA_IN[30]), .CK(net18965), .RN(RST), 
        .Q(\REGISTERS[22][30] ) );
  DFFR_X1 \REGISTERS_reg[22][29]  ( .D(DATA_IN[29]), .CK(net18965), .RN(RST), 
        .Q(\REGISTERS[22][29] ) );
  DFFR_X1 \REGISTERS_reg[22][28]  ( .D(DATA_IN[28]), .CK(net18965), .RN(RST), 
        .Q(\REGISTERS[22][28] ) );
  DFFR_X1 \REGISTERS_reg[22][27]  ( .D(DATA_IN[27]), .CK(net18965), .RN(RST), 
        .Q(\REGISTERS[22][27] ) );
  DFFR_X1 \REGISTERS_reg[22][26]  ( .D(DATA_IN[26]), .CK(net18965), .RN(RST), 
        .Q(\REGISTERS[22][26] ) );
  DFFR_X1 \REGISTERS_reg[22][25]  ( .D(DATA_IN[25]), .CK(net18965), .RN(RST), 
        .Q(\REGISTERS[22][25] ) );
  DFFR_X1 \REGISTERS_reg[22][24]  ( .D(DATA_IN[24]), .CK(net18965), .RN(RST), 
        .Q(\REGISTERS[22][24] ) );
  DFFR_X1 \REGISTERS_reg[22][23]  ( .D(DATA_IN[23]), .CK(net18965), .RN(RST), 
        .Q(\REGISTERS[22][23] ) );
  DFFR_X1 \REGISTERS_reg[22][22]  ( .D(DATA_IN[22]), .CK(net18965), .RN(RST), 
        .Q(\REGISTERS[22][22] ) );
  DFFR_X1 \REGISTERS_reg[22][21]  ( .D(DATA_IN[21]), .CK(net18965), .RN(RST), 
        .Q(\REGISTERS[22][21] ) );
  DFFR_X1 \REGISTERS_reg[22][20]  ( .D(DATA_IN[20]), .CK(net18965), .RN(RST), 
        .Q(\REGISTERS[22][20] ) );
  DFFR_X1 \REGISTERS_reg[22][19]  ( .D(DATA_IN[19]), .CK(net18965), .RN(RST), 
        .Q(\REGISTERS[22][19] ) );
  DFFR_X1 \REGISTERS_reg[22][18]  ( .D(DATA_IN[18]), .CK(net18965), .RN(RST), 
        .Q(\REGISTERS[22][18] ) );
  DFFR_X1 \REGISTERS_reg[22][17]  ( .D(DATA_IN[17]), .CK(net18965), .RN(RST), 
        .Q(\REGISTERS[22][17] ) );
  DFFR_X1 \REGISTERS_reg[22][16]  ( .D(DATA_IN[16]), .CK(net18965), .RN(RST), 
        .Q(\REGISTERS[22][16] ) );
  DFFR_X1 \REGISTERS_reg[22][15]  ( .D(DATA_IN[15]), .CK(net18965), .RN(RST), 
        .Q(\REGISTERS[22][15] ) );
  DFFR_X1 \REGISTERS_reg[22][14]  ( .D(DATA_IN[14]), .CK(net18965), .RN(RST), 
        .Q(\REGISTERS[22][14] ) );
  DFFR_X1 \REGISTERS_reg[22][13]  ( .D(DATA_IN[13]), .CK(net18965), .RN(RST), 
        .Q(\REGISTERS[22][13] ) );
  DFFR_X1 \REGISTERS_reg[22][12]  ( .D(DATA_IN[12]), .CK(net18965), .RN(RST), 
        .Q(\REGISTERS[22][12] ) );
  DFFR_X1 \REGISTERS_reg[22][11]  ( .D(DATA_IN[11]), .CK(net18965), .RN(RST), 
        .Q(\REGISTERS[22][11] ) );
  DFFR_X1 \REGISTERS_reg[22][10]  ( .D(DATA_IN[10]), .CK(net18965), .RN(RST), 
        .Q(\REGISTERS[22][10] ) );
  DFFR_X1 \REGISTERS_reg[22][9]  ( .D(DATA_IN[9]), .CK(net18965), .RN(RST), 
        .Q(\REGISTERS[22][9] ) );
  DFFR_X1 \REGISTERS_reg[22][8]  ( .D(DATA_IN[8]), .CK(net18965), .RN(RST), 
        .Q(\REGISTERS[22][8] ) );
  DFFR_X1 \REGISTERS_reg[22][7]  ( .D(DATA_IN[7]), .CK(net18965), .RN(RST), 
        .Q(\REGISTERS[22][7] ) );
  DFFR_X1 \REGISTERS_reg[22][6]  ( .D(DATA_IN[6]), .CK(net18965), .RN(RST), 
        .Q(\REGISTERS[22][6] ) );
  DFFR_X1 \REGISTERS_reg[22][5]  ( .D(DATA_IN[5]), .CK(net18965), .RN(RST), 
        .Q(\REGISTERS[22][5] ) );
  DFFR_X1 \REGISTERS_reg[22][4]  ( .D(DATA_IN[4]), .CK(net18965), .RN(RST), 
        .Q(\REGISTERS[22][4] ) );
  DFFR_X1 \REGISTERS_reg[22][3]  ( .D(DATA_IN[3]), .CK(net18965), .RN(RST), 
        .Q(\REGISTERS[22][3] ) );
  DFFR_X1 \REGISTERS_reg[22][2]  ( .D(DATA_IN[2]), .CK(net18965), .RN(RST), 
        .Q(\REGISTERS[22][2] ) );
  DFFR_X1 \REGISTERS_reg[22][1]  ( .D(DATA_IN[1]), .CK(net18965), .RN(RST), 
        .Q(\REGISTERS[22][1] ) );
  DFFR_X1 \REGISTERS_reg[22][0]  ( .D(DATA_IN[0]), .CK(net18965), .RN(RST), 
        .Q(\REGISTERS[22][0] ) );
  DFFR_X1 \REGISTERS_reg[23][31]  ( .D(DATA_IN[31]), .CK(net18970), .RN(RST), 
        .Q(\REGISTERS[23][31] ) );
  DFFR_X1 \REGISTERS_reg[23][30]  ( .D(DATA_IN[30]), .CK(net18970), .RN(RST), 
        .Q(\REGISTERS[23][30] ) );
  DFFR_X1 \REGISTERS_reg[23][29]  ( .D(DATA_IN[29]), .CK(net18970), .RN(RST), 
        .Q(\REGISTERS[23][29] ) );
  DFFR_X1 \REGISTERS_reg[23][28]  ( .D(DATA_IN[28]), .CK(net18970), .RN(RST), 
        .Q(\REGISTERS[23][28] ) );
  DFFR_X1 \REGISTERS_reg[23][27]  ( .D(DATA_IN[27]), .CK(net18970), .RN(RST), 
        .Q(\REGISTERS[23][27] ) );
  DFFR_X1 \REGISTERS_reg[23][26]  ( .D(DATA_IN[26]), .CK(net18970), .RN(RST), 
        .Q(\REGISTERS[23][26] ) );
  DFFR_X1 \REGISTERS_reg[23][25]  ( .D(DATA_IN[25]), .CK(net18970), .RN(RST), 
        .Q(\REGISTERS[23][25] ) );
  DFFR_X1 \REGISTERS_reg[23][24]  ( .D(DATA_IN[24]), .CK(net18970), .RN(RST), 
        .Q(\REGISTERS[23][24] ) );
  DFFR_X1 \REGISTERS_reg[23][23]  ( .D(DATA_IN[23]), .CK(net18970), .RN(RST), 
        .Q(\REGISTERS[23][23] ) );
  DFFR_X1 \REGISTERS_reg[23][22]  ( .D(DATA_IN[22]), .CK(net18970), .RN(RST), 
        .Q(\REGISTERS[23][22] ) );
  DFFR_X1 \REGISTERS_reg[23][21]  ( .D(DATA_IN[21]), .CK(net18970), .RN(RST), 
        .Q(\REGISTERS[23][21] ) );
  DFFR_X1 \REGISTERS_reg[23][20]  ( .D(DATA_IN[20]), .CK(net18970), .RN(RST), 
        .Q(\REGISTERS[23][20] ) );
  DFFR_X1 \REGISTERS_reg[23][19]  ( .D(DATA_IN[19]), .CK(net18970), .RN(RST), 
        .Q(\REGISTERS[23][19] ) );
  DFFR_X1 \REGISTERS_reg[23][18]  ( .D(DATA_IN[18]), .CK(net18970), .RN(RST), 
        .Q(\REGISTERS[23][18] ) );
  DFFR_X1 \REGISTERS_reg[23][17]  ( .D(DATA_IN[17]), .CK(net18970), .RN(RST), 
        .Q(\REGISTERS[23][17] ) );
  DFFR_X1 \REGISTERS_reg[23][16]  ( .D(DATA_IN[16]), .CK(net18970), .RN(RST), 
        .Q(\REGISTERS[23][16] ) );
  DFFR_X1 \REGISTERS_reg[23][15]  ( .D(DATA_IN[15]), .CK(net18970), .RN(RST), 
        .Q(\REGISTERS[23][15] ) );
  DFFR_X1 \REGISTERS_reg[23][14]  ( .D(DATA_IN[14]), .CK(net18970), .RN(RST), 
        .Q(\REGISTERS[23][14] ) );
  DFFR_X1 \REGISTERS_reg[23][13]  ( .D(DATA_IN[13]), .CK(net18970), .RN(RST), 
        .Q(\REGISTERS[23][13] ) );
  DFFR_X1 \REGISTERS_reg[23][12]  ( .D(DATA_IN[12]), .CK(net18970), .RN(RST), 
        .Q(\REGISTERS[23][12] ) );
  DFFR_X1 \REGISTERS_reg[23][11]  ( .D(DATA_IN[11]), .CK(net18970), .RN(RST), 
        .Q(\REGISTERS[23][11] ) );
  DFFR_X1 \REGISTERS_reg[23][10]  ( .D(DATA_IN[10]), .CK(net18970), .RN(RST), 
        .Q(\REGISTERS[23][10] ) );
  DFFR_X1 \REGISTERS_reg[23][9]  ( .D(DATA_IN[9]), .CK(net18970), .RN(RST), 
        .Q(\REGISTERS[23][9] ) );
  DFFR_X1 \REGISTERS_reg[23][8]  ( .D(DATA_IN[8]), .CK(net18970), .RN(RST), 
        .Q(\REGISTERS[23][8] ) );
  DFFR_X1 \REGISTERS_reg[23][7]  ( .D(DATA_IN[7]), .CK(net18970), .RN(RST), 
        .Q(\REGISTERS[23][7] ) );
  DFFR_X1 \REGISTERS_reg[23][6]  ( .D(DATA_IN[6]), .CK(net18970), .RN(RST), 
        .Q(\REGISTERS[23][6] ) );
  DFFR_X1 \REGISTERS_reg[23][5]  ( .D(DATA_IN[5]), .CK(net18970), .RN(RST), 
        .Q(\REGISTERS[23][5] ) );
  DFFR_X1 \REGISTERS_reg[23][4]  ( .D(DATA_IN[4]), .CK(net18970), .RN(RST), 
        .Q(\REGISTERS[23][4] ) );
  DFFR_X1 \REGISTERS_reg[23][3]  ( .D(DATA_IN[3]), .CK(net18970), .RN(RST), 
        .Q(\REGISTERS[23][3] ) );
  DFFR_X1 \REGISTERS_reg[23][2]  ( .D(DATA_IN[2]), .CK(net18970), .RN(RST), 
        .Q(\REGISTERS[23][2] ) );
  DFFR_X1 \REGISTERS_reg[23][1]  ( .D(DATA_IN[1]), .CK(net18970), .RN(RST), 
        .Q(\REGISTERS[23][1] ) );
  DFFR_X1 \REGISTERS_reg[23][0]  ( .D(DATA_IN[0]), .CK(net18970), .RN(RST), 
        .Q(\REGISTERS[23][0] ) );
  DFFR_X1 \REGISTERS_reg[24][31]  ( .D(DATA_IN[31]), .CK(net18975), .RN(RST), 
        .Q(\REGISTERS[24][31] ) );
  DFFR_X1 \REGISTERS_reg[24][30]  ( .D(DATA_IN[30]), .CK(net18975), .RN(RST), 
        .Q(\REGISTERS[24][30] ) );
  DFFR_X1 \REGISTERS_reg[24][29]  ( .D(DATA_IN[29]), .CK(net18975), .RN(RST), 
        .Q(\REGISTERS[24][29] ) );
  DFFR_X1 \REGISTERS_reg[24][28]  ( .D(DATA_IN[28]), .CK(net18975), .RN(RST), 
        .Q(\REGISTERS[24][28] ) );
  DFFR_X1 \REGISTERS_reg[24][27]  ( .D(DATA_IN[27]), .CK(net18975), .RN(RST), 
        .Q(\REGISTERS[24][27] ) );
  DFFR_X1 \REGISTERS_reg[24][26]  ( .D(DATA_IN[26]), .CK(net18975), .RN(RST), 
        .Q(\REGISTERS[24][26] ) );
  DFFR_X1 \REGISTERS_reg[24][25]  ( .D(DATA_IN[25]), .CK(net18975), .RN(RST), 
        .Q(\REGISTERS[24][25] ) );
  DFFR_X1 \REGISTERS_reg[24][24]  ( .D(DATA_IN[24]), .CK(net18975), .RN(RST), 
        .Q(\REGISTERS[24][24] ) );
  DFFR_X1 \REGISTERS_reg[24][23]  ( .D(DATA_IN[23]), .CK(net18975), .RN(RST), 
        .Q(\REGISTERS[24][23] ) );
  DFFR_X1 \REGISTERS_reg[24][22]  ( .D(DATA_IN[22]), .CK(net18975), .RN(RST), 
        .Q(\REGISTERS[24][22] ) );
  DFFR_X1 \REGISTERS_reg[24][21]  ( .D(DATA_IN[21]), .CK(net18975), .RN(RST), 
        .Q(\REGISTERS[24][21] ) );
  DFFR_X1 \REGISTERS_reg[24][20]  ( .D(DATA_IN[20]), .CK(net18975), .RN(RST), 
        .Q(\REGISTERS[24][20] ) );
  DFFR_X1 \REGISTERS_reg[24][19]  ( .D(DATA_IN[19]), .CK(net18975), .RN(RST), 
        .Q(\REGISTERS[24][19] ) );
  DFFR_X1 \REGISTERS_reg[24][18]  ( .D(DATA_IN[18]), .CK(net18975), .RN(RST), 
        .Q(\REGISTERS[24][18] ) );
  DFFR_X1 \REGISTERS_reg[24][17]  ( .D(DATA_IN[17]), .CK(net18975), .RN(RST), 
        .Q(\REGISTERS[24][17] ) );
  DFFR_X1 \REGISTERS_reg[24][16]  ( .D(DATA_IN[16]), .CK(net18975), .RN(RST), 
        .Q(\REGISTERS[24][16] ) );
  DFFR_X1 \REGISTERS_reg[24][15]  ( .D(DATA_IN[15]), .CK(net18975), .RN(RST), 
        .Q(\REGISTERS[24][15] ) );
  DFFR_X1 \REGISTERS_reg[24][14]  ( .D(DATA_IN[14]), .CK(net18975), .RN(RST), 
        .Q(\REGISTERS[24][14] ) );
  DFFR_X1 \REGISTERS_reg[24][13]  ( .D(DATA_IN[13]), .CK(net18975), .RN(RST), 
        .Q(\REGISTERS[24][13] ) );
  DFFR_X1 \REGISTERS_reg[24][12]  ( .D(DATA_IN[12]), .CK(net18975), .RN(RST), 
        .Q(\REGISTERS[24][12] ) );
  DFFR_X1 \REGISTERS_reg[24][11]  ( .D(DATA_IN[11]), .CK(net18975), .RN(RST), 
        .Q(\REGISTERS[24][11] ) );
  DFFR_X1 \REGISTERS_reg[24][10]  ( .D(DATA_IN[10]), .CK(net18975), .RN(RST), 
        .Q(\REGISTERS[24][10] ) );
  DFFR_X1 \REGISTERS_reg[24][9]  ( .D(DATA_IN[9]), .CK(net18975), .RN(RST), 
        .Q(\REGISTERS[24][9] ) );
  DFFR_X1 \REGISTERS_reg[24][8]  ( .D(DATA_IN[8]), .CK(net18975), .RN(RST), 
        .Q(\REGISTERS[24][8] ) );
  DFFR_X1 \REGISTERS_reg[24][7]  ( .D(DATA_IN[7]), .CK(net18975), .RN(RST), 
        .Q(\REGISTERS[24][7] ) );
  DFFR_X1 \REGISTERS_reg[24][6]  ( .D(DATA_IN[6]), .CK(net18975), .RN(RST), 
        .Q(\REGISTERS[24][6] ) );
  DFFR_X1 \REGISTERS_reg[24][5]  ( .D(DATA_IN[5]), .CK(net18975), .RN(RST), 
        .Q(\REGISTERS[24][5] ) );
  DFFR_X1 \REGISTERS_reg[24][4]  ( .D(DATA_IN[4]), .CK(net18975), .RN(RST), 
        .Q(\REGISTERS[24][4] ) );
  DFFR_X1 \REGISTERS_reg[24][3]  ( .D(DATA_IN[3]), .CK(net18975), .RN(RST), 
        .Q(\REGISTERS[24][3] ) );
  DFFR_X1 \REGISTERS_reg[24][2]  ( .D(DATA_IN[2]), .CK(net18975), .RN(RST), 
        .Q(\REGISTERS[24][2] ) );
  DFFR_X1 \REGISTERS_reg[24][1]  ( .D(DATA_IN[1]), .CK(net18975), .RN(RST), 
        .Q(\REGISTERS[24][1] ) );
  DFFR_X1 \REGISTERS_reg[24][0]  ( .D(DATA_IN[0]), .CK(net18975), .RN(RST), 
        .Q(\REGISTERS[24][0] ) );
  DFFR_X1 \REGISTERS_reg[25][31]  ( .D(DATA_IN[31]), .CK(net18980), .RN(RST), 
        .Q(\REGISTERS[25][31] ) );
  DFFR_X1 \REGISTERS_reg[25][30]  ( .D(DATA_IN[30]), .CK(net18980), .RN(RST), 
        .Q(\REGISTERS[25][30] ) );
  DFFR_X1 \REGISTERS_reg[25][29]  ( .D(DATA_IN[29]), .CK(net18980), .RN(RST), 
        .Q(\REGISTERS[25][29] ) );
  DFFR_X1 \REGISTERS_reg[25][28]  ( .D(DATA_IN[28]), .CK(net18980), .RN(RST), 
        .Q(\REGISTERS[25][28] ) );
  DFFR_X1 \REGISTERS_reg[25][27]  ( .D(DATA_IN[27]), .CK(net18980), .RN(RST), 
        .Q(\REGISTERS[25][27] ) );
  DFFR_X1 \REGISTERS_reg[25][26]  ( .D(DATA_IN[26]), .CK(net18980), .RN(RST), 
        .Q(\REGISTERS[25][26] ) );
  DFFR_X1 \REGISTERS_reg[25][25]  ( .D(DATA_IN[25]), .CK(net18980), .RN(RST), 
        .Q(\REGISTERS[25][25] ) );
  DFFR_X1 \REGISTERS_reg[25][24]  ( .D(DATA_IN[24]), .CK(net18980), .RN(RST), 
        .Q(\REGISTERS[25][24] ) );
  DFFR_X1 \REGISTERS_reg[25][23]  ( .D(DATA_IN[23]), .CK(net18980), .RN(RST), 
        .Q(\REGISTERS[25][23] ) );
  DFFR_X1 \REGISTERS_reg[25][22]  ( .D(DATA_IN[22]), .CK(net18980), .RN(RST), 
        .Q(\REGISTERS[25][22] ) );
  DFFR_X1 \REGISTERS_reg[25][21]  ( .D(DATA_IN[21]), .CK(net18980), .RN(RST), 
        .Q(\REGISTERS[25][21] ) );
  DFFR_X1 \REGISTERS_reg[25][20]  ( .D(DATA_IN[20]), .CK(net18980), .RN(RST), 
        .Q(\REGISTERS[25][20] ) );
  DFFR_X1 \REGISTERS_reg[25][19]  ( .D(DATA_IN[19]), .CK(net18980), .RN(RST), 
        .Q(\REGISTERS[25][19] ) );
  DFFR_X1 \REGISTERS_reg[25][18]  ( .D(DATA_IN[18]), .CK(net18980), .RN(RST), 
        .Q(\REGISTERS[25][18] ) );
  DFFR_X1 \REGISTERS_reg[25][17]  ( .D(DATA_IN[17]), .CK(net18980), .RN(RST), 
        .Q(\REGISTERS[25][17] ) );
  DFFR_X1 \REGISTERS_reg[25][16]  ( .D(DATA_IN[16]), .CK(net18980), .RN(RST), 
        .Q(\REGISTERS[25][16] ) );
  DFFR_X1 \REGISTERS_reg[25][15]  ( .D(DATA_IN[15]), .CK(net18980), .RN(RST), 
        .Q(\REGISTERS[25][15] ) );
  DFFR_X1 \REGISTERS_reg[25][14]  ( .D(DATA_IN[14]), .CK(net18980), .RN(RST), 
        .Q(\REGISTERS[25][14] ) );
  DFFR_X1 \REGISTERS_reg[25][13]  ( .D(DATA_IN[13]), .CK(net18980), .RN(RST), 
        .Q(\REGISTERS[25][13] ) );
  DFFR_X1 \REGISTERS_reg[25][12]  ( .D(DATA_IN[12]), .CK(net18980), .RN(RST), 
        .Q(\REGISTERS[25][12] ) );
  DFFR_X1 \REGISTERS_reg[25][11]  ( .D(DATA_IN[11]), .CK(net18980), .RN(RST), 
        .Q(\REGISTERS[25][11] ) );
  DFFR_X1 \REGISTERS_reg[25][10]  ( .D(DATA_IN[10]), .CK(net18980), .RN(RST), 
        .Q(\REGISTERS[25][10] ) );
  DFFR_X1 \REGISTERS_reg[25][9]  ( .D(DATA_IN[9]), .CK(net18980), .RN(RST), 
        .Q(\REGISTERS[25][9] ) );
  DFFR_X1 \REGISTERS_reg[25][8]  ( .D(DATA_IN[8]), .CK(net18980), .RN(RST), 
        .Q(\REGISTERS[25][8] ) );
  DFFR_X1 \REGISTERS_reg[25][7]  ( .D(DATA_IN[7]), .CK(net18980), .RN(RST), 
        .Q(\REGISTERS[25][7] ) );
  DFFR_X1 \REGISTERS_reg[25][6]  ( .D(DATA_IN[6]), .CK(net18980), .RN(RST), 
        .Q(\REGISTERS[25][6] ) );
  DFFR_X1 \REGISTERS_reg[25][5]  ( .D(DATA_IN[5]), .CK(net18980), .RN(RST), 
        .Q(\REGISTERS[25][5] ) );
  DFFR_X1 \REGISTERS_reg[25][4]  ( .D(DATA_IN[4]), .CK(net18980), .RN(RST), 
        .Q(\REGISTERS[25][4] ) );
  DFFR_X1 \REGISTERS_reg[25][3]  ( .D(DATA_IN[3]), .CK(net18980), .RN(RST), 
        .Q(\REGISTERS[25][3] ) );
  DFFR_X1 \REGISTERS_reg[25][2]  ( .D(DATA_IN[2]), .CK(net18980), .RN(RST), 
        .Q(\REGISTERS[25][2] ) );
  DFFR_X1 \REGISTERS_reg[25][1]  ( .D(DATA_IN[1]), .CK(net18980), .RN(RST), 
        .Q(\REGISTERS[25][1] ) );
  DFFR_X1 \REGISTERS_reg[25][0]  ( .D(DATA_IN[0]), .CK(net18980), .RN(RST), 
        .Q(\REGISTERS[25][0] ) );
  DFFR_X1 \REGISTERS_reg[26][31]  ( .D(DATA_IN[31]), .CK(net18985), .RN(RST), 
        .Q(\REGISTERS[26][31] ) );
  DFFR_X1 \REGISTERS_reg[26][30]  ( .D(DATA_IN[30]), .CK(net18985), .RN(RST), 
        .Q(\REGISTERS[26][30] ) );
  DFFR_X1 \REGISTERS_reg[26][29]  ( .D(DATA_IN[29]), .CK(net18985), .RN(RST), 
        .Q(\REGISTERS[26][29] ) );
  DFFR_X1 \REGISTERS_reg[26][28]  ( .D(DATA_IN[28]), .CK(net18985), .RN(RST), 
        .Q(\REGISTERS[26][28] ) );
  DFFR_X1 \REGISTERS_reg[26][27]  ( .D(DATA_IN[27]), .CK(net18985), .RN(RST), 
        .Q(\REGISTERS[26][27] ) );
  DFFR_X1 \REGISTERS_reg[26][26]  ( .D(DATA_IN[26]), .CK(net18985), .RN(RST), 
        .Q(\REGISTERS[26][26] ) );
  DFFR_X1 \REGISTERS_reg[26][25]  ( .D(DATA_IN[25]), .CK(net18985), .RN(RST), 
        .Q(\REGISTERS[26][25] ) );
  DFFR_X1 \REGISTERS_reg[26][24]  ( .D(DATA_IN[24]), .CK(net18985), .RN(RST), 
        .Q(\REGISTERS[26][24] ) );
  DFFR_X1 \REGISTERS_reg[26][23]  ( .D(DATA_IN[23]), .CK(net18985), .RN(RST), 
        .Q(\REGISTERS[26][23] ) );
  DFFR_X1 \REGISTERS_reg[26][22]  ( .D(DATA_IN[22]), .CK(net18985), .RN(RST), 
        .Q(\REGISTERS[26][22] ) );
  DFFR_X1 \REGISTERS_reg[26][21]  ( .D(DATA_IN[21]), .CK(net18985), .RN(RST), 
        .Q(\REGISTERS[26][21] ) );
  DFFR_X1 \REGISTERS_reg[26][20]  ( .D(DATA_IN[20]), .CK(net18985), .RN(RST), 
        .Q(\REGISTERS[26][20] ) );
  DFFR_X1 \REGISTERS_reg[26][19]  ( .D(DATA_IN[19]), .CK(net18985), .RN(RST), 
        .Q(\REGISTERS[26][19] ) );
  DFFR_X1 \REGISTERS_reg[26][18]  ( .D(DATA_IN[18]), .CK(net18985), .RN(RST), 
        .Q(\REGISTERS[26][18] ) );
  DFFR_X1 \REGISTERS_reg[26][17]  ( .D(DATA_IN[17]), .CK(net18985), .RN(RST), 
        .Q(\REGISTERS[26][17] ) );
  DFFR_X1 \REGISTERS_reg[26][16]  ( .D(DATA_IN[16]), .CK(net18985), .RN(RST), 
        .Q(\REGISTERS[26][16] ) );
  DFFR_X1 \REGISTERS_reg[26][15]  ( .D(DATA_IN[15]), .CK(net18985), .RN(RST), 
        .Q(\REGISTERS[26][15] ) );
  DFFR_X1 \REGISTERS_reg[26][14]  ( .D(DATA_IN[14]), .CK(net18985), .RN(RST), 
        .Q(\REGISTERS[26][14] ) );
  DFFR_X1 \REGISTERS_reg[26][13]  ( .D(DATA_IN[13]), .CK(net18985), .RN(RST), 
        .Q(\REGISTERS[26][13] ) );
  DFFR_X1 \REGISTERS_reg[26][12]  ( .D(DATA_IN[12]), .CK(net18985), .RN(RST), 
        .Q(\REGISTERS[26][12] ) );
  DFFR_X1 \REGISTERS_reg[26][11]  ( .D(DATA_IN[11]), .CK(net18985), .RN(RST), 
        .Q(\REGISTERS[26][11] ) );
  DFFR_X1 \REGISTERS_reg[26][10]  ( .D(DATA_IN[10]), .CK(net18985), .RN(RST), 
        .Q(\REGISTERS[26][10] ) );
  DFFR_X1 \REGISTERS_reg[26][9]  ( .D(DATA_IN[9]), .CK(net18985), .RN(RST), 
        .Q(\REGISTERS[26][9] ) );
  DFFR_X1 \REGISTERS_reg[26][8]  ( .D(DATA_IN[8]), .CK(net18985), .RN(RST), 
        .Q(\REGISTERS[26][8] ) );
  DFFR_X1 \REGISTERS_reg[26][7]  ( .D(DATA_IN[7]), .CK(net18985), .RN(RST), 
        .Q(\REGISTERS[26][7] ) );
  DFFR_X1 \REGISTERS_reg[26][6]  ( .D(DATA_IN[6]), .CK(net18985), .RN(RST), 
        .Q(\REGISTERS[26][6] ) );
  DFFR_X1 \REGISTERS_reg[26][5]  ( .D(DATA_IN[5]), .CK(net18985), .RN(RST), 
        .Q(\REGISTERS[26][5] ) );
  DFFR_X1 \REGISTERS_reg[26][4]  ( .D(DATA_IN[4]), .CK(net18985), .RN(RST), 
        .Q(\REGISTERS[26][4] ) );
  DFFR_X1 \REGISTERS_reg[26][3]  ( .D(DATA_IN[3]), .CK(net18985), .RN(RST), 
        .Q(\REGISTERS[26][3] ) );
  DFFR_X1 \REGISTERS_reg[26][2]  ( .D(DATA_IN[2]), .CK(net18985), .RN(RST), 
        .Q(\REGISTERS[26][2] ) );
  DFFR_X1 \REGISTERS_reg[26][1]  ( .D(DATA_IN[1]), .CK(net18985), .RN(RST), 
        .Q(\REGISTERS[26][1] ) );
  DFFR_X1 \REGISTERS_reg[26][0]  ( .D(DATA_IN[0]), .CK(net18985), .RN(RST), 
        .Q(\REGISTERS[26][0] ) );
  DFFR_X1 \REGISTERS_reg[27][31]  ( .D(DATA_IN[31]), .CK(net18990), .RN(RST), 
        .Q(\REGISTERS[27][31] ) );
  DFFR_X1 \REGISTERS_reg[27][30]  ( .D(DATA_IN[30]), .CK(net18990), .RN(RST), 
        .Q(\REGISTERS[27][30] ) );
  DFFR_X1 \REGISTERS_reg[27][29]  ( .D(DATA_IN[29]), .CK(net18990), .RN(RST), 
        .Q(\REGISTERS[27][29] ) );
  DFFR_X1 \REGISTERS_reg[27][28]  ( .D(DATA_IN[28]), .CK(net18990), .RN(RST), 
        .Q(\REGISTERS[27][28] ) );
  DFFR_X1 \REGISTERS_reg[27][27]  ( .D(DATA_IN[27]), .CK(net18990), .RN(RST), 
        .Q(\REGISTERS[27][27] ) );
  DFFR_X1 \REGISTERS_reg[27][26]  ( .D(DATA_IN[26]), .CK(net18990), .RN(RST), 
        .Q(\REGISTERS[27][26] ) );
  DFFR_X1 \REGISTERS_reg[27][25]  ( .D(DATA_IN[25]), .CK(net18990), .RN(RST), 
        .Q(\REGISTERS[27][25] ) );
  DFFR_X1 \REGISTERS_reg[27][24]  ( .D(DATA_IN[24]), .CK(net18990), .RN(RST), 
        .Q(\REGISTERS[27][24] ) );
  DFFR_X1 \REGISTERS_reg[27][23]  ( .D(DATA_IN[23]), .CK(net18990), .RN(RST), 
        .Q(\REGISTERS[27][23] ) );
  DFFR_X1 \REGISTERS_reg[27][22]  ( .D(DATA_IN[22]), .CK(net18990), .RN(RST), 
        .Q(\REGISTERS[27][22] ) );
  DFFR_X1 \REGISTERS_reg[27][21]  ( .D(DATA_IN[21]), .CK(net18990), .RN(RST), 
        .Q(\REGISTERS[27][21] ) );
  DFFR_X1 \REGISTERS_reg[27][20]  ( .D(DATA_IN[20]), .CK(net18990), .RN(RST), 
        .Q(\REGISTERS[27][20] ) );
  DFFR_X1 \REGISTERS_reg[27][19]  ( .D(DATA_IN[19]), .CK(net18990), .RN(RST), 
        .Q(\REGISTERS[27][19] ) );
  DFFR_X1 \REGISTERS_reg[27][18]  ( .D(DATA_IN[18]), .CK(net18990), .RN(RST), 
        .Q(\REGISTERS[27][18] ) );
  DFFR_X1 \REGISTERS_reg[27][17]  ( .D(DATA_IN[17]), .CK(net18990), .RN(RST), 
        .Q(\REGISTERS[27][17] ) );
  DFFR_X1 \REGISTERS_reg[27][16]  ( .D(DATA_IN[16]), .CK(net18990), .RN(RST), 
        .Q(\REGISTERS[27][16] ) );
  DFFR_X1 \REGISTERS_reg[27][15]  ( .D(DATA_IN[15]), .CK(net18990), .RN(RST), 
        .Q(\REGISTERS[27][15] ) );
  DFFR_X1 \REGISTERS_reg[27][14]  ( .D(DATA_IN[14]), .CK(net18990), .RN(RST), 
        .Q(\REGISTERS[27][14] ) );
  DFFR_X1 \REGISTERS_reg[27][13]  ( .D(DATA_IN[13]), .CK(net18990), .RN(RST), 
        .Q(\REGISTERS[27][13] ) );
  DFFR_X1 \REGISTERS_reg[27][12]  ( .D(DATA_IN[12]), .CK(net18990), .RN(RST), 
        .Q(\REGISTERS[27][12] ) );
  DFFR_X1 \REGISTERS_reg[27][11]  ( .D(DATA_IN[11]), .CK(net18990), .RN(RST), 
        .Q(\REGISTERS[27][11] ) );
  DFFR_X1 \REGISTERS_reg[27][10]  ( .D(DATA_IN[10]), .CK(net18990), .RN(RST), 
        .Q(\REGISTERS[27][10] ) );
  DFFR_X1 \REGISTERS_reg[27][9]  ( .D(DATA_IN[9]), .CK(net18990), .RN(RST), 
        .Q(\REGISTERS[27][9] ) );
  DFFR_X1 \REGISTERS_reg[27][8]  ( .D(DATA_IN[8]), .CK(net18990), .RN(RST), 
        .Q(\REGISTERS[27][8] ) );
  DFFR_X1 \REGISTERS_reg[27][7]  ( .D(DATA_IN[7]), .CK(net18990), .RN(RST), 
        .Q(\REGISTERS[27][7] ) );
  DFFR_X1 \REGISTERS_reg[27][6]  ( .D(DATA_IN[6]), .CK(net18990), .RN(RST), 
        .Q(\REGISTERS[27][6] ) );
  DFFR_X1 \REGISTERS_reg[27][5]  ( .D(DATA_IN[5]), .CK(net18990), .RN(RST), 
        .Q(\REGISTERS[27][5] ) );
  DFFR_X1 \REGISTERS_reg[27][4]  ( .D(DATA_IN[4]), .CK(net18990), .RN(RST), 
        .Q(\REGISTERS[27][4] ) );
  DFFR_X1 \REGISTERS_reg[27][3]  ( .D(DATA_IN[3]), .CK(net18990), .RN(RST), 
        .Q(\REGISTERS[27][3] ) );
  DFFR_X1 \REGISTERS_reg[27][2]  ( .D(DATA_IN[2]), .CK(net18990), .RN(RST), 
        .Q(\REGISTERS[27][2] ) );
  DFFR_X1 \REGISTERS_reg[27][1]  ( .D(DATA_IN[1]), .CK(net18990), .RN(RST), 
        .Q(\REGISTERS[27][1] ) );
  DFFR_X1 \REGISTERS_reg[27][0]  ( .D(DATA_IN[0]), .CK(net18990), .RN(RST), 
        .Q(\REGISTERS[27][0] ) );
  DFFR_X1 \REGISTERS_reg[28][31]  ( .D(DATA_IN[31]), .CK(net18995), .RN(RST), 
        .Q(\REGISTERS[28][31] ) );
  DFFR_X1 \REGISTERS_reg[28][30]  ( .D(DATA_IN[30]), .CK(net18995), .RN(RST), 
        .Q(\REGISTERS[28][30] ) );
  DFFR_X1 \REGISTERS_reg[28][29]  ( .D(DATA_IN[29]), .CK(net18995), .RN(RST), 
        .Q(\REGISTERS[28][29] ) );
  DFFR_X1 \REGISTERS_reg[28][28]  ( .D(DATA_IN[28]), .CK(net18995), .RN(RST), 
        .Q(\REGISTERS[28][28] ) );
  DFFR_X1 \REGISTERS_reg[28][27]  ( .D(DATA_IN[27]), .CK(net18995), .RN(RST), 
        .Q(\REGISTERS[28][27] ) );
  DFFR_X1 \REGISTERS_reg[28][26]  ( .D(DATA_IN[26]), .CK(net18995), .RN(RST), 
        .Q(\REGISTERS[28][26] ) );
  DFFR_X1 \REGISTERS_reg[28][25]  ( .D(DATA_IN[25]), .CK(net18995), .RN(RST), 
        .Q(\REGISTERS[28][25] ) );
  DFFR_X1 \REGISTERS_reg[28][24]  ( .D(DATA_IN[24]), .CK(net18995), .RN(RST), 
        .Q(\REGISTERS[28][24] ) );
  DFFR_X1 \REGISTERS_reg[28][23]  ( .D(DATA_IN[23]), .CK(net18995), .RN(RST), 
        .Q(\REGISTERS[28][23] ) );
  DFFR_X1 \REGISTERS_reg[28][22]  ( .D(DATA_IN[22]), .CK(net18995), .RN(RST), 
        .Q(\REGISTERS[28][22] ) );
  DFFR_X1 \REGISTERS_reg[28][21]  ( .D(DATA_IN[21]), .CK(net18995), .RN(RST), 
        .Q(\REGISTERS[28][21] ) );
  DFFR_X1 \REGISTERS_reg[28][20]  ( .D(DATA_IN[20]), .CK(net18995), .RN(RST), 
        .Q(\REGISTERS[28][20] ) );
  DFFR_X1 \REGISTERS_reg[28][19]  ( .D(DATA_IN[19]), .CK(net18995), .RN(RST), 
        .Q(\REGISTERS[28][19] ) );
  DFFR_X1 \REGISTERS_reg[28][18]  ( .D(DATA_IN[18]), .CK(net18995), .RN(RST), 
        .Q(\REGISTERS[28][18] ) );
  DFFR_X1 \REGISTERS_reg[28][17]  ( .D(DATA_IN[17]), .CK(net18995), .RN(RST), 
        .Q(\REGISTERS[28][17] ) );
  DFFR_X1 \REGISTERS_reg[28][16]  ( .D(DATA_IN[16]), .CK(net18995), .RN(RST), 
        .Q(\REGISTERS[28][16] ) );
  DFFR_X1 \REGISTERS_reg[28][15]  ( .D(DATA_IN[15]), .CK(net18995), .RN(RST), 
        .Q(\REGISTERS[28][15] ) );
  DFFR_X1 \REGISTERS_reg[28][14]  ( .D(DATA_IN[14]), .CK(net18995), .RN(RST), 
        .Q(\REGISTERS[28][14] ) );
  DFFR_X1 \REGISTERS_reg[28][13]  ( .D(DATA_IN[13]), .CK(net18995), .RN(RST), 
        .Q(\REGISTERS[28][13] ) );
  DFFR_X1 \REGISTERS_reg[28][12]  ( .D(DATA_IN[12]), .CK(net18995), .RN(RST), 
        .Q(\REGISTERS[28][12] ) );
  DFFR_X1 \REGISTERS_reg[28][11]  ( .D(DATA_IN[11]), .CK(net18995), .RN(RST), 
        .Q(\REGISTERS[28][11] ) );
  DFFR_X1 \REGISTERS_reg[28][10]  ( .D(DATA_IN[10]), .CK(net18995), .RN(RST), 
        .Q(\REGISTERS[28][10] ) );
  DFFR_X1 \REGISTERS_reg[28][9]  ( .D(DATA_IN[9]), .CK(net18995), .RN(RST), 
        .Q(\REGISTERS[28][9] ) );
  DFFR_X1 \REGISTERS_reg[28][8]  ( .D(DATA_IN[8]), .CK(net18995), .RN(RST), 
        .Q(\REGISTERS[28][8] ) );
  DFFR_X1 \REGISTERS_reg[28][7]  ( .D(DATA_IN[7]), .CK(net18995), .RN(RST), 
        .Q(\REGISTERS[28][7] ) );
  DFFR_X1 \REGISTERS_reg[28][6]  ( .D(DATA_IN[6]), .CK(net18995), .RN(RST), 
        .Q(\REGISTERS[28][6] ) );
  DFFR_X1 \REGISTERS_reg[28][5]  ( .D(DATA_IN[5]), .CK(net18995), .RN(RST), 
        .Q(\REGISTERS[28][5] ) );
  DFFR_X1 \REGISTERS_reg[28][4]  ( .D(DATA_IN[4]), .CK(net18995), .RN(RST), 
        .Q(\REGISTERS[28][4] ) );
  DFFR_X1 \REGISTERS_reg[28][3]  ( .D(DATA_IN[3]), .CK(net18995), .RN(RST), 
        .Q(\REGISTERS[28][3] ) );
  DFFR_X1 \REGISTERS_reg[28][2]  ( .D(DATA_IN[2]), .CK(net18995), .RN(RST), 
        .Q(\REGISTERS[28][2] ) );
  DFFR_X1 \REGISTERS_reg[28][1]  ( .D(DATA_IN[1]), .CK(net18995), .RN(RST), 
        .Q(\REGISTERS[28][1] ) );
  DFFR_X1 \REGISTERS_reg[28][0]  ( .D(DATA_IN[0]), .CK(net18995), .RN(RST), 
        .Q(\REGISTERS[28][0] ) );
  DFFR_X1 \REGISTERS_reg[29][31]  ( .D(DATA_IN[31]), .CK(net19000), .RN(RST), 
        .Q(\REGISTERS[29][31] ) );
  DFFR_X1 \REGISTERS_reg[29][30]  ( .D(DATA_IN[30]), .CK(net19000), .RN(RST), 
        .Q(\REGISTERS[29][30] ) );
  DFFR_X1 \REGISTERS_reg[29][29]  ( .D(DATA_IN[29]), .CK(net19000), .RN(RST), 
        .Q(\REGISTERS[29][29] ) );
  DFFR_X1 \REGISTERS_reg[29][28]  ( .D(DATA_IN[28]), .CK(net19000), .RN(RST), 
        .Q(\REGISTERS[29][28] ) );
  DFFR_X1 \REGISTERS_reg[29][27]  ( .D(DATA_IN[27]), .CK(net19000), .RN(RST), 
        .Q(\REGISTERS[29][27] ) );
  DFFR_X1 \REGISTERS_reg[29][26]  ( .D(DATA_IN[26]), .CK(net19000), .RN(RST), 
        .Q(\REGISTERS[29][26] ) );
  DFFR_X1 \REGISTERS_reg[29][25]  ( .D(DATA_IN[25]), .CK(net19000), .RN(RST), 
        .Q(\REGISTERS[29][25] ) );
  DFFR_X1 \REGISTERS_reg[29][24]  ( .D(DATA_IN[24]), .CK(net19000), .RN(RST), 
        .Q(\REGISTERS[29][24] ) );
  DFFR_X1 \REGISTERS_reg[29][23]  ( .D(DATA_IN[23]), .CK(net19000), .RN(RST), 
        .Q(\REGISTERS[29][23] ) );
  DFFR_X1 \REGISTERS_reg[29][22]  ( .D(DATA_IN[22]), .CK(net19000), .RN(RST), 
        .Q(\REGISTERS[29][22] ) );
  DFFR_X1 \REGISTERS_reg[29][21]  ( .D(DATA_IN[21]), .CK(net19000), .RN(RST), 
        .Q(\REGISTERS[29][21] ) );
  DFFR_X1 \REGISTERS_reg[29][20]  ( .D(DATA_IN[20]), .CK(net19000), .RN(RST), 
        .Q(\REGISTERS[29][20] ) );
  DFFR_X1 \REGISTERS_reg[29][19]  ( .D(DATA_IN[19]), .CK(net19000), .RN(RST), 
        .Q(\REGISTERS[29][19] ) );
  DFFR_X1 \REGISTERS_reg[29][18]  ( .D(DATA_IN[18]), .CK(net19000), .RN(RST), 
        .Q(\REGISTERS[29][18] ) );
  DFFR_X1 \REGISTERS_reg[29][17]  ( .D(DATA_IN[17]), .CK(net19000), .RN(RST), 
        .Q(\REGISTERS[29][17] ) );
  DFFR_X1 \REGISTERS_reg[29][16]  ( .D(DATA_IN[16]), .CK(net19000), .RN(RST), 
        .Q(\REGISTERS[29][16] ) );
  DFFR_X1 \REGISTERS_reg[29][15]  ( .D(DATA_IN[15]), .CK(net19000), .RN(RST), 
        .Q(\REGISTERS[29][15] ) );
  DFFR_X1 \REGISTERS_reg[29][14]  ( .D(DATA_IN[14]), .CK(net19000), .RN(RST), 
        .Q(\REGISTERS[29][14] ) );
  DFFR_X1 \REGISTERS_reg[29][13]  ( .D(DATA_IN[13]), .CK(net19000), .RN(RST), 
        .Q(\REGISTERS[29][13] ) );
  DFFR_X1 \REGISTERS_reg[29][12]  ( .D(DATA_IN[12]), .CK(net19000), .RN(RST), 
        .Q(\REGISTERS[29][12] ) );
  DFFR_X1 \REGISTERS_reg[29][11]  ( .D(DATA_IN[11]), .CK(net19000), .RN(RST), 
        .Q(\REGISTERS[29][11] ) );
  DFFR_X1 \REGISTERS_reg[29][10]  ( .D(DATA_IN[10]), .CK(net19000), .RN(RST), 
        .Q(\REGISTERS[29][10] ) );
  DFFR_X1 \REGISTERS_reg[29][9]  ( .D(DATA_IN[9]), .CK(net19000), .RN(RST), 
        .Q(\REGISTERS[29][9] ) );
  DFFR_X1 \REGISTERS_reg[29][8]  ( .D(DATA_IN[8]), .CK(net19000), .RN(RST), 
        .Q(\REGISTERS[29][8] ) );
  DFFR_X1 \REGISTERS_reg[29][7]  ( .D(DATA_IN[7]), .CK(net19000), .RN(RST), 
        .Q(\REGISTERS[29][7] ) );
  DFFR_X1 \REGISTERS_reg[29][6]  ( .D(DATA_IN[6]), .CK(net19000), .RN(RST), 
        .Q(\REGISTERS[29][6] ) );
  DFFR_X1 \REGISTERS_reg[29][5]  ( .D(DATA_IN[5]), .CK(net19000), .RN(RST), 
        .Q(\REGISTERS[29][5] ) );
  DFFR_X1 \REGISTERS_reg[29][4]  ( .D(DATA_IN[4]), .CK(net19000), .RN(RST), 
        .Q(\REGISTERS[29][4] ) );
  DFFR_X1 \REGISTERS_reg[29][3]  ( .D(DATA_IN[3]), .CK(net19000), .RN(RST), 
        .Q(\REGISTERS[29][3] ) );
  DFFR_X1 \REGISTERS_reg[29][2]  ( .D(DATA_IN[2]), .CK(net19000), .RN(RST), 
        .Q(\REGISTERS[29][2] ) );
  DFFR_X1 \REGISTERS_reg[29][1]  ( .D(DATA_IN[1]), .CK(net19000), .RN(RST), 
        .Q(\REGISTERS[29][1] ) );
  DFFR_X1 \REGISTERS_reg[29][0]  ( .D(DATA_IN[0]), .CK(net19000), .RN(RST), 
        .Q(\REGISTERS[29][0] ) );
  DFFR_X1 \REGISTERS_reg[30][31]  ( .D(DATA_IN[31]), .CK(net19005), .RN(RST), 
        .Q(\REGISTERS[30][31] ) );
  DFFR_X1 \REGISTERS_reg[30][30]  ( .D(DATA_IN[30]), .CK(net19005), .RN(RST), 
        .Q(\REGISTERS[30][30] ) );
  DFFR_X1 \REGISTERS_reg[30][29]  ( .D(DATA_IN[29]), .CK(net19005), .RN(RST), 
        .Q(\REGISTERS[30][29] ) );
  DFFR_X1 \REGISTERS_reg[30][28]  ( .D(DATA_IN[28]), .CK(net19005), .RN(RST), 
        .Q(\REGISTERS[30][28] ) );
  DFFR_X1 \REGISTERS_reg[30][27]  ( .D(DATA_IN[27]), .CK(net19005), .RN(RST), 
        .Q(\REGISTERS[30][27] ) );
  DFFR_X1 \REGISTERS_reg[30][26]  ( .D(DATA_IN[26]), .CK(net19005), .RN(RST), 
        .Q(\REGISTERS[30][26] ) );
  DFFR_X1 \REGISTERS_reg[30][25]  ( .D(DATA_IN[25]), .CK(net19005), .RN(RST), 
        .Q(\REGISTERS[30][25] ) );
  DFFR_X1 \REGISTERS_reg[30][24]  ( .D(DATA_IN[24]), .CK(net19005), .RN(RST), 
        .Q(\REGISTERS[30][24] ) );
  DFFR_X1 \REGISTERS_reg[30][23]  ( .D(DATA_IN[23]), .CK(net19005), .RN(RST), 
        .Q(\REGISTERS[30][23] ) );
  DFFR_X1 \REGISTERS_reg[30][22]  ( .D(DATA_IN[22]), .CK(net19005), .RN(RST), 
        .Q(\REGISTERS[30][22] ) );
  DFFR_X1 \REGISTERS_reg[30][21]  ( .D(DATA_IN[21]), .CK(net19005), .RN(RST), 
        .Q(\REGISTERS[30][21] ) );
  DFFR_X1 \REGISTERS_reg[30][20]  ( .D(DATA_IN[20]), .CK(net19005), .RN(RST), 
        .Q(\REGISTERS[30][20] ) );
  DFFR_X1 \REGISTERS_reg[30][19]  ( .D(DATA_IN[19]), .CK(net19005), .RN(RST), 
        .Q(\REGISTERS[30][19] ) );
  DFFR_X1 \REGISTERS_reg[30][18]  ( .D(DATA_IN[18]), .CK(net19005), .RN(RST), 
        .Q(\REGISTERS[30][18] ) );
  DFFR_X1 \REGISTERS_reg[30][17]  ( .D(DATA_IN[17]), .CK(net19005), .RN(RST), 
        .Q(\REGISTERS[30][17] ) );
  DFFR_X1 \REGISTERS_reg[30][16]  ( .D(DATA_IN[16]), .CK(net19005), .RN(RST), 
        .Q(\REGISTERS[30][16] ) );
  DFFR_X1 \REGISTERS_reg[30][15]  ( .D(DATA_IN[15]), .CK(net19005), .RN(RST), 
        .Q(\REGISTERS[30][15] ) );
  DFFR_X1 \REGISTERS_reg[30][14]  ( .D(DATA_IN[14]), .CK(net19005), .RN(RST), 
        .Q(\REGISTERS[30][14] ) );
  DFFR_X1 \REGISTERS_reg[30][13]  ( .D(DATA_IN[13]), .CK(net19005), .RN(RST), 
        .Q(\REGISTERS[30][13] ) );
  DFFR_X1 \REGISTERS_reg[30][12]  ( .D(DATA_IN[12]), .CK(net19005), .RN(RST), 
        .Q(\REGISTERS[30][12] ) );
  DFFR_X1 \REGISTERS_reg[30][11]  ( .D(DATA_IN[11]), .CK(net19005), .RN(RST), 
        .Q(\REGISTERS[30][11] ) );
  DFFR_X1 \REGISTERS_reg[30][10]  ( .D(DATA_IN[10]), .CK(net19005), .RN(RST), 
        .Q(\REGISTERS[30][10] ) );
  DFFR_X1 \REGISTERS_reg[30][9]  ( .D(DATA_IN[9]), .CK(net19005), .RN(RST), 
        .Q(\REGISTERS[30][9] ) );
  DFFR_X1 \REGISTERS_reg[30][8]  ( .D(DATA_IN[8]), .CK(net19005), .RN(RST), 
        .Q(\REGISTERS[30][8] ) );
  DFFR_X1 \REGISTERS_reg[30][7]  ( .D(DATA_IN[7]), .CK(net19005), .RN(RST), 
        .Q(\REGISTERS[30][7] ) );
  DFFR_X1 \REGISTERS_reg[30][6]  ( .D(DATA_IN[6]), .CK(net19005), .RN(RST), 
        .Q(\REGISTERS[30][6] ) );
  DFFR_X1 \REGISTERS_reg[30][5]  ( .D(DATA_IN[5]), .CK(net19005), .RN(RST), 
        .Q(\REGISTERS[30][5] ) );
  DFFR_X1 \REGISTERS_reg[30][4]  ( .D(DATA_IN[4]), .CK(net19005), .RN(RST), 
        .Q(\REGISTERS[30][4] ) );
  DFFR_X1 \REGISTERS_reg[30][3]  ( .D(DATA_IN[3]), .CK(net19005), .RN(RST), 
        .Q(\REGISTERS[30][3] ) );
  DFFR_X1 \REGISTERS_reg[30][2]  ( .D(DATA_IN[2]), .CK(net19005), .RN(RST), 
        .Q(\REGISTERS[30][2] ) );
  DFFR_X1 \REGISTERS_reg[30][1]  ( .D(DATA_IN[1]), .CK(net19005), .RN(RST), 
        .Q(\REGISTERS[30][1] ) );
  DFFR_X1 \REGISTERS_reg[30][0]  ( .D(DATA_IN[0]), .CK(net19005), .RN(RST), 
        .Q(\REGISTERS[30][0] ) );
  DFFR_X1 \REGISTERS_reg[31][31]  ( .D(DATA_IN[31]), .CK(net19010), .RN(RST), 
        .Q(\REGISTERS[31][31] ) );
  DFFR_X1 \REGISTERS_reg[31][30]  ( .D(DATA_IN[30]), .CK(net19010), .RN(RST), 
        .Q(\REGISTERS[31][30] ) );
  DFFR_X1 \REGISTERS_reg[31][29]  ( .D(DATA_IN[29]), .CK(net19010), .RN(RST), 
        .Q(\REGISTERS[31][29] ) );
  DFFR_X1 \REGISTERS_reg[31][28]  ( .D(DATA_IN[28]), .CK(net19010), .RN(RST), 
        .Q(\REGISTERS[31][28] ) );
  DFFR_X1 \REGISTERS_reg[31][27]  ( .D(DATA_IN[27]), .CK(net19010), .RN(RST), 
        .Q(\REGISTERS[31][27] ) );
  DFFR_X1 \REGISTERS_reg[31][26]  ( .D(DATA_IN[26]), .CK(net19010), .RN(RST), 
        .Q(\REGISTERS[31][26] ) );
  DFFR_X1 \REGISTERS_reg[31][25]  ( .D(DATA_IN[25]), .CK(net19010), .RN(RST), 
        .Q(\REGISTERS[31][25] ) );
  DFFR_X1 \REGISTERS_reg[31][24]  ( .D(DATA_IN[24]), .CK(net19010), .RN(RST), 
        .Q(\REGISTERS[31][24] ) );
  DFFR_X1 \REGISTERS_reg[31][23]  ( .D(DATA_IN[23]), .CK(net19010), .RN(RST), 
        .Q(\REGISTERS[31][23] ) );
  DFFR_X1 \REGISTERS_reg[31][22]  ( .D(DATA_IN[22]), .CK(net19010), .RN(RST), 
        .Q(\REGISTERS[31][22] ) );
  DFFR_X1 \REGISTERS_reg[31][21]  ( .D(DATA_IN[21]), .CK(net19010), .RN(RST), 
        .Q(\REGISTERS[31][21] ) );
  DFFR_X1 \REGISTERS_reg[31][20]  ( .D(DATA_IN[20]), .CK(net19010), .RN(RST), 
        .Q(\REGISTERS[31][20] ) );
  DFFR_X1 \REGISTERS_reg[31][19]  ( .D(DATA_IN[19]), .CK(net19010), .RN(RST), 
        .Q(\REGISTERS[31][19] ) );
  DFFR_X1 \REGISTERS_reg[31][18]  ( .D(DATA_IN[18]), .CK(net19010), .RN(RST), 
        .Q(\REGISTERS[31][18] ) );
  DFFR_X1 \REGISTERS_reg[31][17]  ( .D(DATA_IN[17]), .CK(net19010), .RN(RST), 
        .Q(\REGISTERS[31][17] ) );
  DFFR_X1 \REGISTERS_reg[31][16]  ( .D(DATA_IN[16]), .CK(net19010), .RN(RST), 
        .Q(\REGISTERS[31][16] ) );
  DFFR_X1 \REGISTERS_reg[31][15]  ( .D(DATA_IN[15]), .CK(net19010), .RN(RST), 
        .Q(\REGISTERS[31][15] ) );
  DFFR_X1 \REGISTERS_reg[31][14]  ( .D(DATA_IN[14]), .CK(net19010), .RN(RST), 
        .Q(\REGISTERS[31][14] ) );
  DFFR_X1 \REGISTERS_reg[31][13]  ( .D(DATA_IN[13]), .CK(net19010), .RN(RST), 
        .Q(\REGISTERS[31][13] ) );
  DFFR_X1 \REGISTERS_reg[31][12]  ( .D(DATA_IN[12]), .CK(net19010), .RN(RST), 
        .Q(\REGISTERS[31][12] ) );
  DFFR_X1 \REGISTERS_reg[31][11]  ( .D(DATA_IN[11]), .CK(net19010), .RN(RST), 
        .Q(\REGISTERS[31][11] ) );
  DFFR_X1 \REGISTERS_reg[31][10]  ( .D(DATA_IN[10]), .CK(net19010), .RN(RST), 
        .Q(\REGISTERS[31][10] ) );
  DFFR_X1 \REGISTERS_reg[31][9]  ( .D(DATA_IN[9]), .CK(net19010), .RN(RST), 
        .Q(\REGISTERS[31][9] ) );
  DFFR_X1 \REGISTERS_reg[31][8]  ( .D(DATA_IN[8]), .CK(net19010), .RN(RST), 
        .Q(\REGISTERS[31][8] ) );
  DFFR_X1 \REGISTERS_reg[31][7]  ( .D(DATA_IN[7]), .CK(net19010), .RN(RST), 
        .Q(\REGISTERS[31][7] ) );
  DFFR_X1 \REGISTERS_reg[31][6]  ( .D(DATA_IN[6]), .CK(net19010), .RN(RST), 
        .Q(\REGISTERS[31][6] ) );
  DFFR_X1 \REGISTERS_reg[31][5]  ( .D(DATA_IN[5]), .CK(net19010), .RN(RST), 
        .Q(\REGISTERS[31][5] ) );
  DFFR_X1 \REGISTERS_reg[31][4]  ( .D(DATA_IN[4]), .CK(net19010), .RN(RST), 
        .Q(\REGISTERS[31][4] ) );
  DFFR_X1 \REGISTERS_reg[31][3]  ( .D(DATA_IN[3]), .CK(net19010), .RN(RST), 
        .Q(\REGISTERS[31][3] ) );
  DFFR_X1 \REGISTERS_reg[31][2]  ( .D(DATA_IN[2]), .CK(net19010), .RN(RST), 
        .Q(\REGISTERS[31][2] ) );
  DFFR_X1 \REGISTERS_reg[31][1]  ( .D(DATA_IN[1]), .CK(net19010), .RN(RST), 
        .Q(\REGISTERS[31][1] ) );
  DFFR_X1 \REGISTERS_reg[31][0]  ( .D(DATA_IN[0]), .CK(net19010), .RN(RST), 
        .Q(\REGISTERS[31][0] ) );
  AOI22_X1 U3 ( .A1(\REGISTERS[19][10] ), .A2(n70), .B1(\REGISTERS[18][10] ), 
        .B2(n71), .ZN(n1) );
  NAND4_X1 U4 ( .A1(n205), .A2(n206), .A3(n1), .A4(n207), .ZN(OUT1[10]) );
  NAND4_X1 U5 ( .A1(n224), .A2(n225), .A3(n226), .A4(n227), .ZN(OUT1[11]) );
  AOI22_X1 U6 ( .A1(\REGISTERS[21][30] ), .A2(n72), .B1(\REGISTERS[20][30] ), 
        .B2(n73), .ZN(n2) );
  AOI22_X1 U7 ( .A1(\REGISTERS[19][30] ), .A2(n70), .B1(\REGISTERS[18][30] ), 
        .B2(n71), .ZN(n3) );
  NAND4_X1 U8 ( .A1(n644), .A2(n645), .A3(n2), .A4(n3), .ZN(OUT1[30]) );
  NAND2_X2 U9 ( .A1(n167), .A2(n166), .ZN(n819) );
  BUF_X1 U10 ( .A(n1486), .Z(n104) );
  BUF_X1 U11 ( .A(n1485), .Z(n103) );
  BUF_X1 U12 ( .A(n790), .Z(n74) );
  BUF_X1 U13 ( .A(n791), .Z(n75) );
  BUF_X1 U14 ( .A(n1484), .Z(n102) );
  BUF_X1 U15 ( .A(n1483), .Z(n101) );
  BUF_X1 U16 ( .A(n1481), .Z(n99) );
  BUF_X1 U17 ( .A(n1482), .Z(n100) );
  BUF_X1 U18 ( .A(n787), .Z(n71) );
  BUF_X1 U19 ( .A(n786), .Z(n70) );
  BUF_X1 U20 ( .A(n789), .Z(n73) );
  BUF_X1 U21 ( .A(n788), .Z(n72) );
  AND2_X2 U22 ( .A1(ADD_RD2[4]), .A2(n867), .ZN(n1520) );
  BUF_X2 U23 ( .A(n1518), .Z(n36) );
  NAND2_X2 U24 ( .A1(n859), .A2(n858), .ZN(n1514) );
  BUF_X2 U25 ( .A(n1519), .Z(n37) );
  NOR4_X2 U26 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[4]), .A3(n177), .A4(n176), .ZN(
        n824) );
  BUF_X1 U27 ( .A(n816), .Z(n92) );
  BUF_X1 U28 ( .A(n817), .Z(n93) );
  BUF_X2 U29 ( .A(n824), .Z(n98) );
  AND2_X2 U30 ( .A1(ADD_RD1[4]), .A2(n175), .ZN(n825) );
  BUF_X2 U31 ( .A(n823), .Z(n97) );
  BUF_X1 U32 ( .A(n822), .Z(n96) );
  BUF_X1 U33 ( .A(n820), .Z(n94) );
  BUF_X1 U34 ( .A(n821), .Z(n95) );
  BUF_X1 U35 ( .A(n810), .Z(n90) );
  BUF_X1 U36 ( .A(n811), .Z(n91) );
  BUF_X1 U37 ( .A(n808), .Z(n88) );
  BUF_X1 U38 ( .A(n809), .Z(n89) );
  BUF_X1 U39 ( .A(n806), .Z(n86) );
  BUF_X1 U40 ( .A(n807), .Z(n87) );
  BUF_X1 U41 ( .A(n804), .Z(n84) );
  BUF_X1 U42 ( .A(n805), .Z(n85) );
  BUF_X1 U43 ( .A(n798), .Z(n82) );
  BUF_X1 U44 ( .A(n799), .Z(n83) );
  BUF_X1 U45 ( .A(n796), .Z(n80) );
  BUF_X1 U46 ( .A(n797), .Z(n81) );
  BUF_X1 U47 ( .A(n794), .Z(n78) );
  BUF_X1 U48 ( .A(n795), .Z(n79) );
  BUF_X1 U49 ( .A(n792), .Z(n76) );
  BUF_X1 U50 ( .A(n793), .Z(n77) );
  NOR2_X1 U51 ( .A1(n174), .A2(n173), .ZN(n822) );
  NOR2_X1 U52 ( .A1(n170), .A2(n176), .ZN(n821) );
  NOR2_X1 U53 ( .A1(n174), .A2(n168), .ZN(n816) );
  NOR2_X1 U54 ( .A1(n176), .A2(n173), .ZN(n810) );
  NOR2_X1 U55 ( .A1(n174), .A2(n161), .ZN(n811) );
  NOR2_X1 U56 ( .A1(n174), .A2(n160), .ZN(n808) );
  NOR2_X1 U57 ( .A1(n159), .A2(n161), .ZN(n809) );
  NOR2_X1 U58 ( .A1(n159), .A2(n160), .ZN(n806) );
  NOR2_X1 U59 ( .A1(n158), .A2(n161), .ZN(n807) );
  NOR2_X1 U60 ( .A1(n158), .A2(n160), .ZN(n804) );
  NOR2_X1 U61 ( .A1(n176), .A2(n161), .ZN(n805) );
  NOR2_X1 U62 ( .A1(n158), .A2(n151), .ZN(n798) );
  NOR2_X1 U63 ( .A1(n159), .A2(n151), .ZN(n799) );
  NOR2_X1 U64 ( .A1(n174), .A2(n151), .ZN(n796) );
  NOR2_X1 U65 ( .A1(n170), .A2(n159), .ZN(n795) );
  NOR2_X1 U66 ( .A1(n158), .A2(n171), .ZN(n792) );
  NOR2_X1 U67 ( .A1(n170), .A2(n158), .ZN(n793) );
  NOR2_X1 U68 ( .A1(ADD_RD1[2]), .A2(n147), .ZN(n790) );
  NOR2_X1 U69 ( .A1(ADD_RD1[1]), .A2(n147), .ZN(n791) );
  NOR2_X1 U70 ( .A1(n159), .A2(n173), .ZN(n788) );
  NOR2_X1 U71 ( .A1(n159), .A2(n168), .ZN(n789) );
  NOR2_X1 U72 ( .A1(n158), .A2(n173), .ZN(n786) );
  NOR2_X1 U73 ( .A1(n158), .A2(n168), .ZN(n787) );
  BUF_X1 U74 ( .A(n1488), .Z(n106) );
  BUF_X1 U75 ( .A(n1490), .Z(n108) );
  BUF_X1 U76 ( .A(n1492), .Z(n110) );
  BUF_X1 U77 ( .A(n1516), .Z(n124) );
  BUF_X1 U78 ( .A(n1512), .Z(n122) );
  BUF_X1 U79 ( .A(n1494), .Z(n112) );
  BUF_X1 U80 ( .A(n1502), .Z(n116) );
  BUF_X1 U81 ( .A(n1504), .Z(n118) );
  BUF_X1 U82 ( .A(n1500), .Z(n114) );
  BUF_X1 U83 ( .A(n1506), .Z(n120) );
  BUF_X1 U84 ( .A(n1489), .Z(n107) );
  BUF_X1 U85 ( .A(n1515), .Z(n123) );
  BUF_X1 U86 ( .A(n1487), .Z(n105) );
  BUF_X1 U87 ( .A(n1493), .Z(n111) );
  BUF_X1 U88 ( .A(n1499), .Z(n113) );
  BUF_X1 U89 ( .A(n1501), .Z(n115) );
  BUF_X1 U90 ( .A(n1505), .Z(n119) );
  BUF_X1 U91 ( .A(n1517), .Z(n125) );
  BUF_X1 U92 ( .A(n1511), .Z(n121) );
  BUF_X1 U93 ( .A(n1491), .Z(n109) );
  BUF_X1 U94 ( .A(n1503), .Z(n117) );
  NAND3_X1 U95 ( .A1(ADD_WR[1]), .A2(ADD_WR[2]), .A3(ADD_WR[0]), .ZN(n137) );
  NAND3_X1 U96 ( .A1(ADD_WR[4]), .A2(ADD_WR[3]), .A3(WR_EN), .ZN(n130) );
  NOR2_X1 U97 ( .A1(n137), .A2(n130), .ZN(N409) );
  INV_X1 U98 ( .A(ADD_WR[0]), .ZN(n126) );
  NAND3_X1 U99 ( .A1(ADD_WR[2]), .A2(ADD_WR[1]), .A3(n126), .ZN(n138) );
  NOR2_X1 U100 ( .A1(n130), .A2(n138), .ZN(N410) );
  INV_X1 U101 ( .A(ADD_WR[1]), .ZN(n128) );
  NAND3_X1 U102 ( .A1(ADD_WR[2]), .A2(ADD_WR[0]), .A3(n128), .ZN(n139) );
  NOR2_X1 U103 ( .A1(n130), .A2(n139), .ZN(N411) );
  NAND3_X1 U104 ( .A1(ADD_WR[2]), .A2(n128), .A3(n126), .ZN(n140) );
  NOR2_X1 U105 ( .A1(n130), .A2(n140), .ZN(N412) );
  NOR2_X1 U106 ( .A1(ADD_WR[2]), .A2(n126), .ZN(n127) );
  NAND2_X1 U107 ( .A1(ADD_WR[1]), .A2(n127), .ZN(n141) );
  NOR2_X1 U108 ( .A1(n130), .A2(n141), .ZN(N413) );
  NOR2_X1 U109 ( .A1(ADD_WR[2]), .A2(ADD_WR[0]), .ZN(n129) );
  NAND2_X1 U110 ( .A1(ADD_WR[1]), .A2(n129), .ZN(n142) );
  NOR2_X1 U111 ( .A1(n130), .A2(n142), .ZN(N414) );
  NAND2_X1 U112 ( .A1(n127), .A2(n128), .ZN(n144) );
  NOR2_X1 U113 ( .A1(n130), .A2(n144), .ZN(N415) );
  NAND2_X1 U114 ( .A1(n129), .A2(n128), .ZN(n134) );
  NOR2_X1 U115 ( .A1(n130), .A2(n134), .ZN(N416) );
  INV_X1 U116 ( .A(WR_EN), .ZN(n131) );
  NOR2_X1 U117 ( .A1(ADD_WR[3]), .A2(n131), .ZN(n136) );
  NAND2_X1 U118 ( .A1(ADD_WR[4]), .A2(n136), .ZN(n132) );
  NOR2_X1 U119 ( .A1(n137), .A2(n132), .ZN(N417) );
  NOR2_X1 U120 ( .A1(n138), .A2(n132), .ZN(N418) );
  NOR2_X1 U121 ( .A1(n139), .A2(n132), .ZN(N419) );
  NOR2_X1 U122 ( .A1(n140), .A2(n132), .ZN(N420) );
  NOR2_X1 U123 ( .A1(n141), .A2(n132), .ZN(N421) );
  NOR2_X1 U124 ( .A1(n142), .A2(n132), .ZN(N422) );
  NOR2_X1 U125 ( .A1(n144), .A2(n132), .ZN(N423) );
  NOR2_X1 U126 ( .A1(n134), .A2(n132), .ZN(N424) );
  INV_X1 U127 ( .A(ADD_WR[4]), .ZN(n135) );
  NAND3_X1 U128 ( .A1(ADD_WR[3]), .A2(WR_EN), .A3(n135), .ZN(n133) );
  NOR2_X1 U129 ( .A1(n137), .A2(n133), .ZN(N425) );
  NOR2_X1 U130 ( .A1(n138), .A2(n133), .ZN(N426) );
  NOR2_X1 U131 ( .A1(n139), .A2(n133), .ZN(N427) );
  NOR2_X1 U132 ( .A1(n140), .A2(n133), .ZN(N428) );
  NOR2_X1 U133 ( .A1(n141), .A2(n133), .ZN(N429) );
  NOR2_X1 U134 ( .A1(n142), .A2(n133), .ZN(N430) );
  NOR2_X1 U135 ( .A1(n144), .A2(n133), .ZN(N431) );
  NOR2_X1 U136 ( .A1(n134), .A2(n133), .ZN(N432) );
  NAND2_X1 U137 ( .A1(n136), .A2(n135), .ZN(n143) );
  NOR2_X1 U138 ( .A1(n137), .A2(n143), .ZN(N433) );
  NOR2_X1 U139 ( .A1(n138), .A2(n143), .ZN(N434) );
  NOR2_X1 U140 ( .A1(n139), .A2(n143), .ZN(N435) );
  NOR2_X1 U141 ( .A1(n140), .A2(n143), .ZN(N436) );
  NOR2_X1 U142 ( .A1(n141), .A2(n143), .ZN(N437) );
  NOR2_X1 U143 ( .A1(n142), .A2(n143), .ZN(N438) );
  NOR2_X1 U144 ( .A1(n144), .A2(n143), .ZN(N439) );
  INV_X1 U145 ( .A(ADD_RD1[2]), .ZN(n148) );
  NAND2_X1 U146 ( .A1(ADD_RD1[1]), .A2(n148), .ZN(n158) );
  INV_X1 U147 ( .A(ADD_RD1[0]), .ZN(n177) );
  INV_X1 U148 ( .A(ADD_RD1[3]), .ZN(n145) );
  NAND3_X1 U149 ( .A1(ADD_RD1[4]), .A2(n177), .A3(n145), .ZN(n168) );
  NAND3_X1 U150 ( .A1(ADD_RD1[4]), .A2(ADD_RD1[0]), .A3(n145), .ZN(n173) );
  AOI22_X1 U151 ( .A1(\REGISTERS[18][0] ), .A2(n71), .B1(\REGISTERS[19][0] ), 
        .B2(n70), .ZN(n188) );
  INV_X1 U152 ( .A(ADD_RD1[1]), .ZN(n149) );
  NAND2_X1 U153 ( .A1(ADD_RD1[2]), .A2(n149), .ZN(n159) );
  AOI22_X1 U154 ( .A1(\REGISTERS[20][0] ), .A2(n73), .B1(\REGISTERS[21][0] ), 
        .B2(n72), .ZN(n187) );
  NOR3_X1 U155 ( .A1(ADD_RD1[0]), .A2(ADD_RD1[4]), .A3(ADD_RD1[3]), .ZN(n166)
         );
  NAND2_X1 U156 ( .A1(n149), .A2(n148), .ZN(n176) );
  NOR3_X1 U157 ( .A1(ADD_RD1[0]), .A2(ADD_RD1[3]), .A3(n176), .ZN(n175) );
  INV_X1 U158 ( .A(ADD_RD1[4]), .ZN(n156) );
  NAND2_X1 U159 ( .A1(n175), .A2(n156), .ZN(n146) );
  NAND2_X1 U160 ( .A1(n166), .A2(n146), .ZN(n147) );
  AOI22_X1 U161 ( .A1(\REGISTERS[4][0] ), .A2(n75), .B1(\REGISTERS[2][0] ), 
        .B2(n74), .ZN(n186) );
  NAND3_X1 U162 ( .A1(ADD_RD1[4]), .A2(ADD_RD1[3]), .A3(n177), .ZN(n170) );
  NAND3_X1 U163 ( .A1(ADD_RD1[0]), .A2(ADD_RD1[4]), .A3(ADD_RD1[3]), .ZN(n171)
         );
  AOI22_X1 U164 ( .A1(\REGISTERS[26][0] ), .A2(n77), .B1(\REGISTERS[27][0] ), 
        .B2(n76), .ZN(n155) );
  NOR2_X1 U165 ( .A1(n171), .A2(n159), .ZN(n794) );
  AOI22_X1 U166 ( .A1(\REGISTERS[28][0] ), .A2(n79), .B1(\REGISTERS[29][0] ), 
        .B2(n78), .ZN(n154) );
  NOR2_X1 U167 ( .A1(n149), .A2(n148), .ZN(n167) );
  INV_X1 U168 ( .A(n167), .ZN(n174) );
  NOR2_X1 U169 ( .A1(n170), .A2(n174), .ZN(n797) );
  NOR2_X1 U170 ( .A1(ADD_RD1[4]), .A2(ADD_RD1[3]), .ZN(n150) );
  NAND2_X1 U171 ( .A1(ADD_RD1[0]), .A2(n150), .ZN(n151) );
  AOI22_X1 U172 ( .A1(\REGISTERS[30][0] ), .A2(n81), .B1(\REGISTERS[7][0] ), 
        .B2(n80), .ZN(n153) );
  AOI22_X1 U173 ( .A1(\REGISTERS[5][0] ), .A2(n83), .B1(\REGISTERS[3][0] ), 
        .B2(n82), .ZN(n152) );
  NAND4_X1 U174 ( .A1(n155), .A2(n154), .A3(n153), .A4(n152), .ZN(n184) );
  NAND2_X1 U175 ( .A1(n156), .A2(ADD_RD1[3]), .ZN(n172) );
  INV_X1 U176 ( .A(n172), .ZN(n157) );
  NAND2_X1 U177 ( .A1(ADD_RD1[0]), .A2(n157), .ZN(n161) );
  NAND2_X1 U178 ( .A1(n157), .A2(n177), .ZN(n160) );
  AOI22_X1 U179 ( .A1(\REGISTERS[9][0] ), .A2(n85), .B1(\REGISTERS[10][0] ), 
        .B2(n84), .ZN(n165) );
  AOI22_X1 U180 ( .A1(\REGISTERS[11][0] ), .A2(n87), .B1(\REGISTERS[12][0] ), 
        .B2(n86), .ZN(n164) );
  AOI22_X1 U181 ( .A1(\REGISTERS[13][0] ), .A2(n89), .B1(\REGISTERS[14][0] ), 
        .B2(n88), .ZN(n163) );
  AOI22_X1 U182 ( .A1(\REGISTERS[15][0] ), .A2(n91), .B1(\REGISTERS[17][0] ), 
        .B2(n90), .ZN(n162) );
  NAND4_X1 U183 ( .A1(n165), .A2(n164), .A3(n163), .A4(n162), .ZN(n183) );
  NOR2_X1 U184 ( .A1(n171), .A2(n174), .ZN(n817) );
  AOI22_X1 U185 ( .A1(\REGISTERS[31][0] ), .A2(n93), .B1(\REGISTERS[22][0] ), 
        .B2(n92), .ZN(n169) );
  OAI21_X1 U186 ( .B1(n38), .B2(n819), .A(n169), .ZN(n182) );
  NOR2_X1 U187 ( .A1(n171), .A2(n176), .ZN(n820) );
  AOI22_X1 U188 ( .A1(\REGISTERS[24][0] ), .A2(n95), .B1(\REGISTERS[25][0] ), 
        .B2(n94), .ZN(n180) );
  NOR3_X1 U189 ( .A1(ADD_RD1[0]), .A2(n176), .A3(n172), .ZN(n823) );
  AOI22_X1 U190 ( .A1(\REGISTERS[8][0] ), .A2(n97), .B1(\REGISTERS[23][0] ), 
        .B2(n96), .ZN(n179) );
  AOI22_X1 U191 ( .A1(\REGISTERS[16][0] ), .A2(n825), .B1(\REGISTERS[1][0] ), 
        .B2(n98), .ZN(n178) );
  NAND3_X1 U192 ( .A1(n180), .A2(n179), .A3(n178), .ZN(n181) );
  NOR4_X1 U193 ( .A1(n184), .A2(n183), .A3(n182), .A4(n181), .ZN(n185) );
  NAND4_X1 U194 ( .A1(n188), .A2(n187), .A3(n186), .A4(n185), .ZN(OUT1[0]) );
  AOI22_X1 U195 ( .A1(n73), .A2(\REGISTERS[20][10] ), .B1(n72), .B2(
        \REGISTERS[21][10] ), .ZN(n207) );
  AOI22_X1 U196 ( .A1(n75), .A2(\REGISTERS[4][10] ), .B1(n74), .B2(
        \REGISTERS[2][10] ), .ZN(n206) );
  AOI22_X1 U197 ( .A1(n77), .A2(\REGISTERS[26][10] ), .B1(n76), .B2(
        \REGISTERS[27][10] ), .ZN(n192) );
  AOI22_X1 U198 ( .A1(n79), .A2(\REGISTERS[28][10] ), .B1(n78), .B2(
        \REGISTERS[29][10] ), .ZN(n191) );
  AOI22_X1 U199 ( .A1(n81), .A2(\REGISTERS[30][10] ), .B1(n80), .B2(
        \REGISTERS[7][10] ), .ZN(n190) );
  AOI22_X1 U200 ( .A1(n83), .A2(\REGISTERS[5][10] ), .B1(n82), .B2(
        \REGISTERS[3][10] ), .ZN(n189) );
  NAND4_X1 U201 ( .A1(n192), .A2(n191), .A3(n190), .A4(n189), .ZN(n204) );
  AOI22_X1 U202 ( .A1(n85), .A2(\REGISTERS[9][10] ), .B1(n84), .B2(
        \REGISTERS[10][10] ), .ZN(n196) );
  AOI22_X1 U203 ( .A1(n87), .A2(\REGISTERS[11][10] ), .B1(n86), .B2(
        \REGISTERS[12][10] ), .ZN(n195) );
  AOI22_X1 U204 ( .A1(n89), .A2(\REGISTERS[13][10] ), .B1(n88), .B2(
        \REGISTERS[14][10] ), .ZN(n194) );
  AOI22_X1 U205 ( .A1(n91), .A2(\REGISTERS[15][10] ), .B1(n90), .B2(
        \REGISTERS[17][10] ), .ZN(n193) );
  NAND4_X1 U206 ( .A1(n196), .A2(n195), .A3(n194), .A4(n193), .ZN(n203) );
  AOI22_X1 U207 ( .A1(n93), .A2(\REGISTERS[31][10] ), .B1(n92), .B2(
        \REGISTERS[22][10] ), .ZN(n197) );
  OAI21_X1 U208 ( .B1(n819), .B2(n39), .A(n197), .ZN(n202) );
  AOI22_X1 U209 ( .A1(n95), .A2(\REGISTERS[24][10] ), .B1(n94), .B2(
        \REGISTERS[25][10] ), .ZN(n200) );
  AOI22_X1 U210 ( .A1(n97), .A2(\REGISTERS[8][10] ), .B1(n96), .B2(
        \REGISTERS[23][10] ), .ZN(n199) );
  AOI22_X1 U211 ( .A1(n825), .A2(\REGISTERS[16][10] ), .B1(n98), .B2(
        \REGISTERS[1][10] ), .ZN(n198) );
  NAND3_X1 U212 ( .A1(n200), .A2(n199), .A3(n198), .ZN(n201) );
  NOR4_X1 U213 ( .A1(n204), .A2(n203), .A3(n202), .A4(n201), .ZN(n205) );
  AOI22_X1 U214 ( .A1(n787), .A2(\REGISTERS[18][11] ), .B1(n786), .B2(
        \REGISTERS[19][11] ), .ZN(n227) );
  AOI22_X1 U215 ( .A1(n789), .A2(\REGISTERS[20][11] ), .B1(n788), .B2(
        \REGISTERS[21][11] ), .ZN(n226) );
  AOI22_X1 U216 ( .A1(n75), .A2(\REGISTERS[4][11] ), .B1(n790), .B2(
        \REGISTERS[2][11] ), .ZN(n225) );
  AOI22_X1 U217 ( .A1(n793), .A2(\REGISTERS[26][11] ), .B1(n792), .B2(
        \REGISTERS[27][11] ), .ZN(n211) );
  AOI22_X1 U218 ( .A1(n795), .A2(\REGISTERS[28][11] ), .B1(n794), .B2(
        \REGISTERS[29][11] ), .ZN(n210) );
  AOI22_X1 U219 ( .A1(n797), .A2(\REGISTERS[30][11] ), .B1(n796), .B2(
        \REGISTERS[7][11] ), .ZN(n209) );
  AOI22_X1 U220 ( .A1(n83), .A2(\REGISTERS[5][11] ), .B1(n798), .B2(
        \REGISTERS[3][11] ), .ZN(n208) );
  NAND4_X1 U221 ( .A1(n211), .A2(n210), .A3(n209), .A4(n208), .ZN(n223) );
  AOI22_X1 U222 ( .A1(n85), .A2(\REGISTERS[9][11] ), .B1(n84), .B2(
        \REGISTERS[10][11] ), .ZN(n215) );
  AOI22_X1 U223 ( .A1(n807), .A2(\REGISTERS[11][11] ), .B1(n86), .B2(
        \REGISTERS[12][11] ), .ZN(n214) );
  AOI22_X1 U224 ( .A1(n809), .A2(\REGISTERS[13][11] ), .B1(n88), .B2(
        \REGISTERS[14][11] ), .ZN(n213) );
  AOI22_X1 U225 ( .A1(n91), .A2(\REGISTERS[15][11] ), .B1(n810), .B2(
        \REGISTERS[17][11] ), .ZN(n212) );
  NAND4_X1 U226 ( .A1(n215), .A2(n214), .A3(n213), .A4(n212), .ZN(n222) );
  AOI22_X1 U227 ( .A1(n817), .A2(\REGISTERS[31][11] ), .B1(n816), .B2(
        \REGISTERS[22][11] ), .ZN(n216) );
  OAI21_X1 U228 ( .B1(n819), .B2(n40), .A(n216), .ZN(n221) );
  AOI22_X1 U229 ( .A1(n821), .A2(\REGISTERS[24][11] ), .B1(n820), .B2(
        \REGISTERS[25][11] ), .ZN(n219) );
  AOI22_X1 U230 ( .A1(n823), .A2(\REGISTERS[8][11] ), .B1(n822), .B2(
        \REGISTERS[23][11] ), .ZN(n218) );
  AOI22_X1 U231 ( .A1(n825), .A2(\REGISTERS[16][11] ), .B1(n98), .B2(
        \REGISTERS[1][11] ), .ZN(n217) );
  NAND3_X1 U232 ( .A1(n219), .A2(n218), .A3(n217), .ZN(n220) );
  NOR4_X1 U233 ( .A1(n223), .A2(n222), .A3(n221), .A4(n220), .ZN(n224) );
  AOI22_X1 U234 ( .A1(n787), .A2(\REGISTERS[18][12] ), .B1(n786), .B2(
        \REGISTERS[19][12] ), .ZN(n247) );
  AOI22_X1 U235 ( .A1(n789), .A2(\REGISTERS[20][12] ), .B1(n788), .B2(
        \REGISTERS[21][12] ), .ZN(n246) );
  AOI22_X1 U236 ( .A1(n75), .A2(\REGISTERS[4][12] ), .B1(n790), .B2(
        \REGISTERS[2][12] ), .ZN(n245) );
  AOI22_X1 U237 ( .A1(n77), .A2(\REGISTERS[26][12] ), .B1(n792), .B2(
        \REGISTERS[27][12] ), .ZN(n231) );
  AOI22_X1 U238 ( .A1(n79), .A2(\REGISTERS[28][12] ), .B1(n794), .B2(
        \REGISTERS[29][12] ), .ZN(n230) );
  AOI22_X1 U239 ( .A1(n81), .A2(\REGISTERS[30][12] ), .B1(n80), .B2(
        \REGISTERS[7][12] ), .ZN(n229) );
  AOI22_X1 U240 ( .A1(n83), .A2(\REGISTERS[5][12] ), .B1(n798), .B2(
        \REGISTERS[3][12] ), .ZN(n228) );
  NAND4_X1 U241 ( .A1(n231), .A2(n230), .A3(n229), .A4(n228), .ZN(n243) );
  AOI22_X1 U242 ( .A1(n85), .A2(\REGISTERS[9][12] ), .B1(n84), .B2(
        \REGISTERS[10][12] ), .ZN(n235) );
  AOI22_X1 U243 ( .A1(n87), .A2(\REGISTERS[11][12] ), .B1(n86), .B2(
        \REGISTERS[12][12] ), .ZN(n234) );
  AOI22_X1 U244 ( .A1(n89), .A2(\REGISTERS[13][12] ), .B1(n88), .B2(
        \REGISTERS[14][12] ), .ZN(n233) );
  AOI22_X1 U245 ( .A1(n91), .A2(\REGISTERS[15][12] ), .B1(n90), .B2(
        \REGISTERS[17][12] ), .ZN(n232) );
  NAND4_X1 U246 ( .A1(n235), .A2(n234), .A3(n233), .A4(n232), .ZN(n242) );
  AOI22_X1 U247 ( .A1(n93), .A2(\REGISTERS[31][12] ), .B1(n92), .B2(
        \REGISTERS[22][12] ), .ZN(n236) );
  OAI21_X1 U248 ( .B1(n819), .B2(n41), .A(n236), .ZN(n241) );
  AOI22_X1 U249 ( .A1(n95), .A2(\REGISTERS[24][12] ), .B1(n94), .B2(
        \REGISTERS[25][12] ), .ZN(n239) );
  AOI22_X1 U250 ( .A1(n97), .A2(\REGISTERS[8][12] ), .B1(n96), .B2(
        \REGISTERS[23][12] ), .ZN(n238) );
  AOI22_X1 U251 ( .A1(n825), .A2(\REGISTERS[16][12] ), .B1(n824), .B2(
        \REGISTERS[1][12] ), .ZN(n237) );
  NAND3_X1 U252 ( .A1(n239), .A2(n238), .A3(n237), .ZN(n240) );
  NOR4_X1 U253 ( .A1(n243), .A2(n242), .A3(n241), .A4(n240), .ZN(n244) );
  NAND4_X1 U254 ( .A1(n247), .A2(n246), .A3(n245), .A4(n244), .ZN(OUT1[12]) );
  AOI22_X1 U255 ( .A1(n71), .A2(\REGISTERS[18][13] ), .B1(n70), .B2(
        \REGISTERS[19][13] ), .ZN(n267) );
  AOI22_X1 U256 ( .A1(n73), .A2(\REGISTERS[20][13] ), .B1(n72), .B2(
        \REGISTERS[21][13] ), .ZN(n266) );
  AOI22_X1 U257 ( .A1(n75), .A2(\REGISTERS[4][13] ), .B1(n74), .B2(
        \REGISTERS[2][13] ), .ZN(n265) );
  AOI22_X1 U258 ( .A1(n77), .A2(\REGISTERS[26][13] ), .B1(n76), .B2(
        \REGISTERS[27][13] ), .ZN(n251) );
  AOI22_X1 U259 ( .A1(n79), .A2(\REGISTERS[28][13] ), .B1(n78), .B2(
        \REGISTERS[29][13] ), .ZN(n250) );
  AOI22_X1 U260 ( .A1(n81), .A2(\REGISTERS[30][13] ), .B1(n80), .B2(
        \REGISTERS[7][13] ), .ZN(n249) );
  AOI22_X1 U261 ( .A1(n83), .A2(\REGISTERS[5][13] ), .B1(n82), .B2(
        \REGISTERS[3][13] ), .ZN(n248) );
  NAND4_X1 U262 ( .A1(n251), .A2(n250), .A3(n249), .A4(n248), .ZN(n263) );
  AOI22_X1 U263 ( .A1(n85), .A2(\REGISTERS[9][13] ), .B1(n84), .B2(
        \REGISTERS[10][13] ), .ZN(n255) );
  AOI22_X1 U264 ( .A1(n87), .A2(\REGISTERS[11][13] ), .B1(n86), .B2(
        \REGISTERS[12][13] ), .ZN(n254) );
  AOI22_X1 U265 ( .A1(n89), .A2(\REGISTERS[13][13] ), .B1(n88), .B2(
        \REGISTERS[14][13] ), .ZN(n253) );
  AOI22_X1 U266 ( .A1(n91), .A2(\REGISTERS[15][13] ), .B1(n90), .B2(
        \REGISTERS[17][13] ), .ZN(n252) );
  NAND4_X1 U267 ( .A1(n255), .A2(n254), .A3(n253), .A4(n252), .ZN(n262) );
  AOI22_X1 U268 ( .A1(n93), .A2(\REGISTERS[31][13] ), .B1(n92), .B2(
        \REGISTERS[22][13] ), .ZN(n256) );
  OAI21_X1 U269 ( .B1(n819), .B2(n42), .A(n256), .ZN(n261) );
  AOI22_X1 U270 ( .A1(n95), .A2(\REGISTERS[24][13] ), .B1(n94), .B2(
        \REGISTERS[25][13] ), .ZN(n259) );
  AOI22_X1 U271 ( .A1(n97), .A2(\REGISTERS[8][13] ), .B1(n96), .B2(
        \REGISTERS[23][13] ), .ZN(n258) );
  AOI22_X1 U272 ( .A1(n825), .A2(\REGISTERS[16][13] ), .B1(n98), .B2(
        \REGISTERS[1][13] ), .ZN(n257) );
  NAND3_X1 U273 ( .A1(n259), .A2(n258), .A3(n257), .ZN(n260) );
  NOR4_X1 U274 ( .A1(n263), .A2(n262), .A3(n261), .A4(n260), .ZN(n264) );
  NAND4_X1 U275 ( .A1(n267), .A2(n266), .A3(n265), .A4(n264), .ZN(OUT1[13]) );
  AOI22_X1 U276 ( .A1(n71), .A2(\REGISTERS[18][14] ), .B1(n70), .B2(
        \REGISTERS[19][14] ), .ZN(n287) );
  AOI22_X1 U277 ( .A1(n73), .A2(\REGISTERS[20][14] ), .B1(n72), .B2(
        \REGISTERS[21][14] ), .ZN(n286) );
  AOI22_X1 U278 ( .A1(n75), .A2(\REGISTERS[4][14] ), .B1(n74), .B2(
        \REGISTERS[2][14] ), .ZN(n285) );
  AOI22_X1 U279 ( .A1(n77), .A2(\REGISTERS[26][14] ), .B1(n76), .B2(
        \REGISTERS[27][14] ), .ZN(n271) );
  AOI22_X1 U280 ( .A1(n79), .A2(\REGISTERS[28][14] ), .B1(n78), .B2(
        \REGISTERS[29][14] ), .ZN(n270) );
  AOI22_X1 U281 ( .A1(n81), .A2(\REGISTERS[30][14] ), .B1(n80), .B2(
        \REGISTERS[7][14] ), .ZN(n269) );
  AOI22_X1 U282 ( .A1(n83), .A2(\REGISTERS[5][14] ), .B1(n82), .B2(
        \REGISTERS[3][14] ), .ZN(n268) );
  NAND4_X1 U283 ( .A1(n271), .A2(n270), .A3(n269), .A4(n268), .ZN(n283) );
  AOI22_X1 U284 ( .A1(n85), .A2(\REGISTERS[9][14] ), .B1(n84), .B2(
        \REGISTERS[10][14] ), .ZN(n275) );
  AOI22_X1 U285 ( .A1(n87), .A2(\REGISTERS[11][14] ), .B1(n86), .B2(
        \REGISTERS[12][14] ), .ZN(n274) );
  AOI22_X1 U286 ( .A1(n89), .A2(\REGISTERS[13][14] ), .B1(n88), .B2(
        \REGISTERS[14][14] ), .ZN(n273) );
  AOI22_X1 U287 ( .A1(n91), .A2(\REGISTERS[15][14] ), .B1(n90), .B2(
        \REGISTERS[17][14] ), .ZN(n272) );
  NAND4_X1 U288 ( .A1(n275), .A2(n274), .A3(n273), .A4(n272), .ZN(n282) );
  AOI22_X1 U289 ( .A1(n93), .A2(\REGISTERS[31][14] ), .B1(n92), .B2(
        \REGISTERS[22][14] ), .ZN(n276) );
  OAI21_X1 U290 ( .B1(n819), .B2(n43), .A(n276), .ZN(n281) );
  AOI22_X1 U291 ( .A1(n95), .A2(\REGISTERS[24][14] ), .B1(n94), .B2(
        \REGISTERS[25][14] ), .ZN(n279) );
  AOI22_X1 U292 ( .A1(n97), .A2(\REGISTERS[8][14] ), .B1(n96), .B2(
        \REGISTERS[23][14] ), .ZN(n278) );
  AOI22_X1 U293 ( .A1(n825), .A2(\REGISTERS[16][14] ), .B1(n98), .B2(
        \REGISTERS[1][14] ), .ZN(n277) );
  NAND3_X1 U294 ( .A1(n279), .A2(n278), .A3(n277), .ZN(n280) );
  NOR4_X1 U295 ( .A1(n283), .A2(n282), .A3(n281), .A4(n280), .ZN(n284) );
  NAND4_X1 U296 ( .A1(n287), .A2(n286), .A3(n285), .A4(n284), .ZN(OUT1[14]) );
  AOI22_X1 U297 ( .A1(n787), .A2(\REGISTERS[18][15] ), .B1(n786), .B2(
        \REGISTERS[19][15] ), .ZN(n307) );
  AOI22_X1 U298 ( .A1(n73), .A2(\REGISTERS[20][15] ), .B1(n788), .B2(
        \REGISTERS[21][15] ), .ZN(n306) );
  AOI22_X1 U299 ( .A1(n791), .A2(\REGISTERS[4][15] ), .B1(n74), .B2(
        \REGISTERS[2][15] ), .ZN(n305) );
  AOI22_X1 U300 ( .A1(n793), .A2(\REGISTERS[26][15] ), .B1(n792), .B2(
        \REGISTERS[27][15] ), .ZN(n291) );
  AOI22_X1 U301 ( .A1(n795), .A2(\REGISTERS[28][15] ), .B1(n794), .B2(
        \REGISTERS[29][15] ), .ZN(n290) );
  AOI22_X1 U302 ( .A1(n797), .A2(\REGISTERS[30][15] ), .B1(n796), .B2(
        \REGISTERS[7][15] ), .ZN(n289) );
  AOI22_X1 U303 ( .A1(n799), .A2(\REGISTERS[5][15] ), .B1(n82), .B2(
        \REGISTERS[3][15] ), .ZN(n288) );
  NAND4_X1 U304 ( .A1(n291), .A2(n290), .A3(n289), .A4(n288), .ZN(n303) );
  AOI22_X1 U305 ( .A1(n805), .A2(\REGISTERS[9][15] ), .B1(n804), .B2(
        \REGISTERS[10][15] ), .ZN(n295) );
  AOI22_X1 U306 ( .A1(n807), .A2(\REGISTERS[11][15] ), .B1(n806), .B2(
        \REGISTERS[12][15] ), .ZN(n294) );
  AOI22_X1 U307 ( .A1(n809), .A2(\REGISTERS[13][15] ), .B1(n808), .B2(
        \REGISTERS[14][15] ), .ZN(n293) );
  AOI22_X1 U308 ( .A1(n811), .A2(\REGISTERS[15][15] ), .B1(n810), .B2(
        \REGISTERS[17][15] ), .ZN(n292) );
  NAND4_X1 U309 ( .A1(n295), .A2(n294), .A3(n293), .A4(n292), .ZN(n302) );
  AOI22_X1 U310 ( .A1(n817), .A2(\REGISTERS[31][15] ), .B1(n816), .B2(
        \REGISTERS[22][15] ), .ZN(n296) );
  OAI21_X1 U311 ( .B1(n819), .B2(n44), .A(n296), .ZN(n301) );
  AOI22_X1 U312 ( .A1(n821), .A2(\REGISTERS[24][15] ), .B1(n820), .B2(
        \REGISTERS[25][15] ), .ZN(n299) );
  AOI22_X1 U313 ( .A1(n97), .A2(\REGISTERS[8][15] ), .B1(n822), .B2(
        \REGISTERS[23][15] ), .ZN(n298) );
  AOI22_X1 U314 ( .A1(n825), .A2(\REGISTERS[16][15] ), .B1(n98), .B2(
        \REGISTERS[1][15] ), .ZN(n297) );
  NAND3_X1 U315 ( .A1(n299), .A2(n298), .A3(n297), .ZN(n300) );
  NOR4_X1 U316 ( .A1(n303), .A2(n302), .A3(n301), .A4(n300), .ZN(n304) );
  NAND4_X1 U317 ( .A1(n307), .A2(n306), .A3(n305), .A4(n304), .ZN(OUT1[15]) );
  AOI22_X1 U318 ( .A1(n787), .A2(\REGISTERS[18][16] ), .B1(n786), .B2(
        \REGISTERS[19][16] ), .ZN(n327) );
  AOI22_X1 U319 ( .A1(n789), .A2(\REGISTERS[20][16] ), .B1(n788), .B2(
        \REGISTERS[21][16] ), .ZN(n326) );
  AOI22_X1 U320 ( .A1(n791), .A2(\REGISTERS[4][16] ), .B1(n790), .B2(
        \REGISTERS[2][16] ), .ZN(n325) );
  AOI22_X1 U321 ( .A1(n793), .A2(\REGISTERS[26][16] ), .B1(n792), .B2(
        \REGISTERS[27][16] ), .ZN(n311) );
  AOI22_X1 U322 ( .A1(n795), .A2(\REGISTERS[28][16] ), .B1(n794), .B2(
        \REGISTERS[29][16] ), .ZN(n310) );
  AOI22_X1 U323 ( .A1(n797), .A2(\REGISTERS[30][16] ), .B1(n796), .B2(
        \REGISTERS[7][16] ), .ZN(n309) );
  AOI22_X1 U324 ( .A1(n799), .A2(\REGISTERS[5][16] ), .B1(n798), .B2(
        \REGISTERS[3][16] ), .ZN(n308) );
  NAND4_X1 U325 ( .A1(n311), .A2(n310), .A3(n309), .A4(n308), .ZN(n323) );
  AOI22_X1 U326 ( .A1(n805), .A2(\REGISTERS[9][16] ), .B1(n804), .B2(
        \REGISTERS[10][16] ), .ZN(n315) );
  AOI22_X1 U327 ( .A1(n807), .A2(\REGISTERS[11][16] ), .B1(n806), .B2(
        \REGISTERS[12][16] ), .ZN(n314) );
  AOI22_X1 U328 ( .A1(n809), .A2(\REGISTERS[13][16] ), .B1(n808), .B2(
        \REGISTERS[14][16] ), .ZN(n313) );
  AOI22_X1 U329 ( .A1(n811), .A2(\REGISTERS[15][16] ), .B1(n810), .B2(
        \REGISTERS[17][16] ), .ZN(n312) );
  NAND4_X1 U330 ( .A1(n315), .A2(n314), .A3(n313), .A4(n312), .ZN(n322) );
  AOI22_X1 U331 ( .A1(n817), .A2(\REGISTERS[31][16] ), .B1(n816), .B2(
        \REGISTERS[22][16] ), .ZN(n316) );
  OAI21_X1 U332 ( .B1(n819), .B2(n45), .A(n316), .ZN(n321) );
  AOI22_X1 U333 ( .A1(n821), .A2(\REGISTERS[24][16] ), .B1(n820), .B2(
        \REGISTERS[25][16] ), .ZN(n319) );
  AOI22_X1 U334 ( .A1(n97), .A2(\REGISTERS[8][16] ), .B1(n822), .B2(
        \REGISTERS[23][16] ), .ZN(n318) );
  AOI22_X1 U335 ( .A1(n825), .A2(\REGISTERS[16][16] ), .B1(n98), .B2(
        \REGISTERS[1][16] ), .ZN(n317) );
  NAND3_X1 U336 ( .A1(n319), .A2(n318), .A3(n317), .ZN(n320) );
  NOR4_X1 U337 ( .A1(n323), .A2(n322), .A3(n321), .A4(n320), .ZN(n324) );
  NAND4_X1 U338 ( .A1(n327), .A2(n326), .A3(n325), .A4(n324), .ZN(OUT1[16]) );
  AOI22_X1 U339 ( .A1(n787), .A2(\REGISTERS[18][17] ), .B1(n786), .B2(
        \REGISTERS[19][17] ), .ZN(n347) );
  AOI22_X1 U340 ( .A1(n789), .A2(\REGISTERS[20][17] ), .B1(n788), .B2(
        \REGISTERS[21][17] ), .ZN(n346) );
  AOI22_X1 U341 ( .A1(n791), .A2(\REGISTERS[4][17] ), .B1(n790), .B2(
        \REGISTERS[2][17] ), .ZN(n345) );
  AOI22_X1 U342 ( .A1(n793), .A2(\REGISTERS[26][17] ), .B1(n792), .B2(
        \REGISTERS[27][17] ), .ZN(n331) );
  AOI22_X1 U343 ( .A1(n795), .A2(\REGISTERS[28][17] ), .B1(n794), .B2(
        \REGISTERS[29][17] ), .ZN(n330) );
  AOI22_X1 U344 ( .A1(n797), .A2(\REGISTERS[30][17] ), .B1(n796), .B2(
        \REGISTERS[7][17] ), .ZN(n329) );
  AOI22_X1 U345 ( .A1(n799), .A2(\REGISTERS[5][17] ), .B1(n798), .B2(
        \REGISTERS[3][17] ), .ZN(n328) );
  NAND4_X1 U346 ( .A1(n331), .A2(n330), .A3(n329), .A4(n328), .ZN(n343) );
  AOI22_X1 U347 ( .A1(n805), .A2(\REGISTERS[9][17] ), .B1(n804), .B2(
        \REGISTERS[10][17] ), .ZN(n335) );
  AOI22_X1 U348 ( .A1(n807), .A2(\REGISTERS[11][17] ), .B1(n806), .B2(
        \REGISTERS[12][17] ), .ZN(n334) );
  AOI22_X1 U349 ( .A1(n809), .A2(\REGISTERS[13][17] ), .B1(n808), .B2(
        \REGISTERS[14][17] ), .ZN(n333) );
  AOI22_X1 U350 ( .A1(n811), .A2(\REGISTERS[15][17] ), .B1(n810), .B2(
        \REGISTERS[17][17] ), .ZN(n332) );
  NAND4_X1 U351 ( .A1(n335), .A2(n334), .A3(n333), .A4(n332), .ZN(n342) );
  AOI22_X1 U352 ( .A1(n817), .A2(\REGISTERS[31][17] ), .B1(n816), .B2(
        \REGISTERS[22][17] ), .ZN(n336) );
  OAI21_X1 U353 ( .B1(n819), .B2(n46), .A(n336), .ZN(n341) );
  AOI22_X1 U354 ( .A1(n821), .A2(\REGISTERS[24][17] ), .B1(n820), .B2(
        \REGISTERS[25][17] ), .ZN(n339) );
  AOI22_X1 U355 ( .A1(n97), .A2(\REGISTERS[8][17] ), .B1(n822), .B2(
        \REGISTERS[23][17] ), .ZN(n338) );
  AOI22_X1 U356 ( .A1(n825), .A2(\REGISTERS[16][17] ), .B1(n98), .B2(
        \REGISTERS[1][17] ), .ZN(n337) );
  NAND3_X1 U357 ( .A1(n339), .A2(n338), .A3(n337), .ZN(n340) );
  NOR4_X1 U358 ( .A1(n343), .A2(n342), .A3(n341), .A4(n340), .ZN(n344) );
  NAND4_X1 U359 ( .A1(n347), .A2(n346), .A3(n345), .A4(n344), .ZN(OUT1[17]) );
  AOI22_X1 U360 ( .A1(n787), .A2(\REGISTERS[18][18] ), .B1(n786), .B2(
        \REGISTERS[19][18] ), .ZN(n367) );
  AOI22_X1 U361 ( .A1(n789), .A2(\REGISTERS[20][18] ), .B1(n788), .B2(
        \REGISTERS[21][18] ), .ZN(n366) );
  AOI22_X1 U362 ( .A1(n791), .A2(\REGISTERS[4][18] ), .B1(n790), .B2(
        \REGISTERS[2][18] ), .ZN(n365) );
  AOI22_X1 U363 ( .A1(n793), .A2(\REGISTERS[26][18] ), .B1(n792), .B2(
        \REGISTERS[27][18] ), .ZN(n351) );
  AOI22_X1 U364 ( .A1(n795), .A2(\REGISTERS[28][18] ), .B1(n794), .B2(
        \REGISTERS[29][18] ), .ZN(n350) );
  AOI22_X1 U365 ( .A1(n81), .A2(\REGISTERS[30][18] ), .B1(n80), .B2(
        \REGISTERS[7][18] ), .ZN(n349) );
  AOI22_X1 U366 ( .A1(n799), .A2(\REGISTERS[5][18] ), .B1(n798), .B2(
        \REGISTERS[3][18] ), .ZN(n348) );
  NAND4_X1 U367 ( .A1(n351), .A2(n350), .A3(n349), .A4(n348), .ZN(n363) );
  AOI22_X1 U368 ( .A1(n805), .A2(\REGISTERS[9][18] ), .B1(n804), .B2(
        \REGISTERS[10][18] ), .ZN(n355) );
  AOI22_X1 U369 ( .A1(n807), .A2(\REGISTERS[11][18] ), .B1(n806), .B2(
        \REGISTERS[12][18] ), .ZN(n354) );
  AOI22_X1 U370 ( .A1(n809), .A2(\REGISTERS[13][18] ), .B1(n808), .B2(
        \REGISTERS[14][18] ), .ZN(n353) );
  AOI22_X1 U371 ( .A1(n811), .A2(\REGISTERS[15][18] ), .B1(n90), .B2(
        \REGISTERS[17][18] ), .ZN(n352) );
  NAND4_X1 U372 ( .A1(n355), .A2(n354), .A3(n353), .A4(n352), .ZN(n362) );
  AOI22_X1 U373 ( .A1(n93), .A2(\REGISTERS[31][18] ), .B1(n92), .B2(
        \REGISTERS[22][18] ), .ZN(n356) );
  OAI21_X1 U374 ( .B1(n819), .B2(n47), .A(n356), .ZN(n361) );
  AOI22_X1 U375 ( .A1(n821), .A2(\REGISTERS[24][18] ), .B1(n94), .B2(
        \REGISTERS[25][18] ), .ZN(n359) );
  AOI22_X1 U376 ( .A1(n97), .A2(\REGISTERS[8][18] ), .B1(n822), .B2(
        \REGISTERS[23][18] ), .ZN(n358) );
  AOI22_X1 U377 ( .A1(n825), .A2(\REGISTERS[16][18] ), .B1(n98), .B2(
        \REGISTERS[1][18] ), .ZN(n357) );
  NAND3_X1 U378 ( .A1(n359), .A2(n358), .A3(n357), .ZN(n360) );
  NOR4_X1 U379 ( .A1(n363), .A2(n362), .A3(n361), .A4(n360), .ZN(n364) );
  NAND4_X1 U380 ( .A1(n367), .A2(n366), .A3(n365), .A4(n364), .ZN(OUT1[18]) );
  AOI22_X1 U381 ( .A1(n71), .A2(\REGISTERS[18][19] ), .B1(n70), .B2(
        \REGISTERS[19][19] ), .ZN(n387) );
  AOI22_X1 U382 ( .A1(n73), .A2(\REGISTERS[20][19] ), .B1(n72), .B2(
        \REGISTERS[21][19] ), .ZN(n386) );
  AOI22_X1 U383 ( .A1(n75), .A2(\REGISTERS[4][19] ), .B1(n74), .B2(
        \REGISTERS[2][19] ), .ZN(n385) );
  AOI22_X1 U384 ( .A1(n77), .A2(\REGISTERS[26][19] ), .B1(n76), .B2(
        \REGISTERS[27][19] ), .ZN(n371) );
  AOI22_X1 U385 ( .A1(n79), .A2(\REGISTERS[28][19] ), .B1(n78), .B2(
        \REGISTERS[29][19] ), .ZN(n370) );
  AOI22_X1 U386 ( .A1(n81), .A2(\REGISTERS[30][19] ), .B1(n80), .B2(
        \REGISTERS[7][19] ), .ZN(n369) );
  AOI22_X1 U387 ( .A1(n83), .A2(\REGISTERS[5][19] ), .B1(n82), .B2(
        \REGISTERS[3][19] ), .ZN(n368) );
  NAND4_X1 U388 ( .A1(n371), .A2(n370), .A3(n369), .A4(n368), .ZN(n383) );
  AOI22_X1 U389 ( .A1(n85), .A2(\REGISTERS[9][19] ), .B1(n84), .B2(
        \REGISTERS[10][19] ), .ZN(n375) );
  AOI22_X1 U390 ( .A1(n87), .A2(\REGISTERS[11][19] ), .B1(n86), .B2(
        \REGISTERS[12][19] ), .ZN(n374) );
  AOI22_X1 U391 ( .A1(n89), .A2(\REGISTERS[13][19] ), .B1(n88), .B2(
        \REGISTERS[14][19] ), .ZN(n373) );
  AOI22_X1 U392 ( .A1(n91), .A2(\REGISTERS[15][19] ), .B1(n90), .B2(
        \REGISTERS[17][19] ), .ZN(n372) );
  NAND4_X1 U393 ( .A1(n375), .A2(n374), .A3(n373), .A4(n372), .ZN(n382) );
  AOI22_X1 U394 ( .A1(n93), .A2(\REGISTERS[31][19] ), .B1(n92), .B2(
        \REGISTERS[22][19] ), .ZN(n376) );
  OAI21_X1 U395 ( .B1(n819), .B2(n48), .A(n376), .ZN(n381) );
  AOI22_X1 U396 ( .A1(n95), .A2(\REGISTERS[24][19] ), .B1(n94), .B2(
        \REGISTERS[25][19] ), .ZN(n379) );
  AOI22_X1 U397 ( .A1(n97), .A2(\REGISTERS[8][19] ), .B1(n96), .B2(
        \REGISTERS[23][19] ), .ZN(n378) );
  AOI22_X1 U398 ( .A1(n825), .A2(\REGISTERS[16][19] ), .B1(n98), .B2(
        \REGISTERS[1][19] ), .ZN(n377) );
  NAND3_X1 U399 ( .A1(n379), .A2(n378), .A3(n377), .ZN(n380) );
  NOR4_X1 U400 ( .A1(n383), .A2(n382), .A3(n381), .A4(n380), .ZN(n384) );
  NAND4_X1 U401 ( .A1(n387), .A2(n386), .A3(n385), .A4(n384), .ZN(OUT1[19]) );
  AOI22_X1 U402 ( .A1(n787), .A2(\REGISTERS[18][1] ), .B1(n786), .B2(
        \REGISTERS[19][1] ), .ZN(n407) );
  AOI22_X1 U403 ( .A1(n789), .A2(\REGISTERS[20][1] ), .B1(n788), .B2(
        \REGISTERS[21][1] ), .ZN(n406) );
  AOI22_X1 U404 ( .A1(n791), .A2(\REGISTERS[4][1] ), .B1(n790), .B2(
        \REGISTERS[2][1] ), .ZN(n405) );
  AOI22_X1 U405 ( .A1(n793), .A2(\REGISTERS[26][1] ), .B1(n792), .B2(
        \REGISTERS[27][1] ), .ZN(n391) );
  AOI22_X1 U406 ( .A1(n795), .A2(\REGISTERS[28][1] ), .B1(n794), .B2(
        \REGISTERS[29][1] ), .ZN(n390) );
  AOI22_X1 U407 ( .A1(n797), .A2(\REGISTERS[30][1] ), .B1(n796), .B2(
        \REGISTERS[7][1] ), .ZN(n389) );
  AOI22_X1 U408 ( .A1(n799), .A2(\REGISTERS[5][1] ), .B1(n798), .B2(
        \REGISTERS[3][1] ), .ZN(n388) );
  NAND4_X1 U409 ( .A1(n391), .A2(n390), .A3(n389), .A4(n388), .ZN(n403) );
  AOI22_X1 U410 ( .A1(n805), .A2(\REGISTERS[9][1] ), .B1(n804), .B2(
        \REGISTERS[10][1] ), .ZN(n395) );
  AOI22_X1 U411 ( .A1(n807), .A2(\REGISTERS[11][1] ), .B1(n806), .B2(
        \REGISTERS[12][1] ), .ZN(n394) );
  AOI22_X1 U412 ( .A1(n809), .A2(\REGISTERS[13][1] ), .B1(n808), .B2(
        \REGISTERS[14][1] ), .ZN(n393) );
  AOI22_X1 U413 ( .A1(n811), .A2(\REGISTERS[15][1] ), .B1(n810), .B2(
        \REGISTERS[17][1] ), .ZN(n392) );
  NAND4_X1 U414 ( .A1(n395), .A2(n394), .A3(n393), .A4(n392), .ZN(n402) );
  AOI22_X1 U415 ( .A1(n817), .A2(\REGISTERS[31][1] ), .B1(n816), .B2(
        \REGISTERS[22][1] ), .ZN(n396) );
  OAI21_X1 U416 ( .B1(n819), .B2(n49), .A(n396), .ZN(n401) );
  AOI22_X1 U417 ( .A1(n821), .A2(\REGISTERS[24][1] ), .B1(n820), .B2(
        \REGISTERS[25][1] ), .ZN(n399) );
  AOI22_X1 U418 ( .A1(n823), .A2(\REGISTERS[8][1] ), .B1(n822), .B2(
        \REGISTERS[23][1] ), .ZN(n398) );
  AOI22_X1 U419 ( .A1(n825), .A2(\REGISTERS[16][1] ), .B1(n824), .B2(
        \REGISTERS[1][1] ), .ZN(n397) );
  NAND3_X1 U420 ( .A1(n399), .A2(n398), .A3(n397), .ZN(n400) );
  NOR4_X1 U421 ( .A1(n403), .A2(n402), .A3(n401), .A4(n400), .ZN(n404) );
  NAND4_X1 U422 ( .A1(n407), .A2(n406), .A3(n405), .A4(n404), .ZN(OUT1[1]) );
  AOI22_X1 U423 ( .A1(n787), .A2(\REGISTERS[18][20] ), .B1(n786), .B2(
        \REGISTERS[19][20] ), .ZN(n427) );
  AOI22_X1 U424 ( .A1(n789), .A2(\REGISTERS[20][20] ), .B1(n788), .B2(
        \REGISTERS[21][20] ), .ZN(n426) );
  AOI22_X1 U425 ( .A1(n791), .A2(\REGISTERS[4][20] ), .B1(n790), .B2(
        \REGISTERS[2][20] ), .ZN(n425) );
  AOI22_X1 U426 ( .A1(n793), .A2(\REGISTERS[26][20] ), .B1(n76), .B2(
        \REGISTERS[27][20] ), .ZN(n411) );
  AOI22_X1 U427 ( .A1(n795), .A2(\REGISTERS[28][20] ), .B1(n794), .B2(
        \REGISTERS[29][20] ), .ZN(n410) );
  AOI22_X1 U428 ( .A1(n797), .A2(\REGISTERS[30][20] ), .B1(n796), .B2(
        \REGISTERS[7][20] ), .ZN(n409) );
  AOI22_X1 U429 ( .A1(n799), .A2(\REGISTERS[5][20] ), .B1(n798), .B2(
        \REGISTERS[3][20] ), .ZN(n408) );
  NAND4_X1 U430 ( .A1(n411), .A2(n410), .A3(n409), .A4(n408), .ZN(n423) );
  AOI22_X1 U431 ( .A1(n805), .A2(\REGISTERS[9][20] ), .B1(n804), .B2(
        \REGISTERS[10][20] ), .ZN(n415) );
  AOI22_X1 U432 ( .A1(n807), .A2(\REGISTERS[11][20] ), .B1(n806), .B2(
        \REGISTERS[12][20] ), .ZN(n414) );
  AOI22_X1 U433 ( .A1(n809), .A2(\REGISTERS[13][20] ), .B1(n808), .B2(
        \REGISTERS[14][20] ), .ZN(n413) );
  AOI22_X1 U434 ( .A1(n811), .A2(\REGISTERS[15][20] ), .B1(n810), .B2(
        \REGISTERS[17][20] ), .ZN(n412) );
  NAND4_X1 U435 ( .A1(n415), .A2(n414), .A3(n413), .A4(n412), .ZN(n422) );
  AOI22_X1 U436 ( .A1(n817), .A2(\REGISTERS[31][20] ), .B1(n816), .B2(
        \REGISTERS[22][20] ), .ZN(n416) );
  OAI21_X1 U437 ( .B1(n819), .B2(n50), .A(n416), .ZN(n421) );
  AOI22_X1 U438 ( .A1(n821), .A2(\REGISTERS[24][20] ), .B1(n820), .B2(
        \REGISTERS[25][20] ), .ZN(n419) );
  AOI22_X1 U439 ( .A1(n823), .A2(\REGISTERS[8][20] ), .B1(n96), .B2(
        \REGISTERS[23][20] ), .ZN(n418) );
  AOI22_X1 U440 ( .A1(n825), .A2(\REGISTERS[16][20] ), .B1(n824), .B2(
        \REGISTERS[1][20] ), .ZN(n417) );
  NAND3_X1 U441 ( .A1(n419), .A2(n418), .A3(n417), .ZN(n420) );
  NOR4_X1 U442 ( .A1(n423), .A2(n422), .A3(n421), .A4(n420), .ZN(n424) );
  NAND4_X1 U443 ( .A1(n427), .A2(n426), .A3(n425), .A4(n424), .ZN(OUT1[20]) );
  AOI22_X1 U444 ( .A1(n71), .A2(\REGISTERS[18][21] ), .B1(n70), .B2(
        \REGISTERS[19][21] ), .ZN(n447) );
  AOI22_X1 U445 ( .A1(n73), .A2(\REGISTERS[20][21] ), .B1(n72), .B2(
        \REGISTERS[21][21] ), .ZN(n446) );
  AOI22_X1 U446 ( .A1(n75), .A2(\REGISTERS[4][21] ), .B1(n74), .B2(
        \REGISTERS[2][21] ), .ZN(n445) );
  AOI22_X1 U447 ( .A1(n77), .A2(\REGISTERS[26][21] ), .B1(n76), .B2(
        \REGISTERS[27][21] ), .ZN(n431) );
  AOI22_X1 U448 ( .A1(n79), .A2(\REGISTERS[28][21] ), .B1(n78), .B2(
        \REGISTERS[29][21] ), .ZN(n430) );
  AOI22_X1 U449 ( .A1(n81), .A2(\REGISTERS[30][21] ), .B1(n80), .B2(
        \REGISTERS[7][21] ), .ZN(n429) );
  AOI22_X1 U450 ( .A1(n83), .A2(\REGISTERS[5][21] ), .B1(n82), .B2(
        \REGISTERS[3][21] ), .ZN(n428) );
  NAND4_X1 U451 ( .A1(n431), .A2(n430), .A3(n429), .A4(n428), .ZN(n443) );
  AOI22_X1 U452 ( .A1(n85), .A2(\REGISTERS[9][21] ), .B1(n84), .B2(
        \REGISTERS[10][21] ), .ZN(n435) );
  AOI22_X1 U453 ( .A1(n87), .A2(\REGISTERS[11][21] ), .B1(n86), .B2(
        \REGISTERS[12][21] ), .ZN(n434) );
  AOI22_X1 U454 ( .A1(n89), .A2(\REGISTERS[13][21] ), .B1(n88), .B2(
        \REGISTERS[14][21] ), .ZN(n433) );
  AOI22_X1 U455 ( .A1(n91), .A2(\REGISTERS[15][21] ), .B1(n90), .B2(
        \REGISTERS[17][21] ), .ZN(n432) );
  NAND4_X1 U456 ( .A1(n435), .A2(n434), .A3(n433), .A4(n432), .ZN(n442) );
  AOI22_X1 U457 ( .A1(n93), .A2(\REGISTERS[31][21] ), .B1(n92), .B2(
        \REGISTERS[22][21] ), .ZN(n436) );
  OAI21_X1 U458 ( .B1(n819), .B2(n51), .A(n436), .ZN(n441) );
  AOI22_X1 U459 ( .A1(n95), .A2(\REGISTERS[24][21] ), .B1(n94), .B2(
        \REGISTERS[25][21] ), .ZN(n439) );
  AOI22_X1 U460 ( .A1(n97), .A2(\REGISTERS[8][21] ), .B1(n96), .B2(
        \REGISTERS[23][21] ), .ZN(n438) );
  AOI22_X1 U461 ( .A1(n825), .A2(\REGISTERS[16][21] ), .B1(n98), .B2(
        \REGISTERS[1][21] ), .ZN(n437) );
  NAND3_X1 U462 ( .A1(n439), .A2(n438), .A3(n437), .ZN(n440) );
  NOR4_X1 U463 ( .A1(n443), .A2(n442), .A3(n441), .A4(n440), .ZN(n444) );
  NAND4_X1 U464 ( .A1(n447), .A2(n446), .A3(n445), .A4(n444), .ZN(OUT1[21]) );
  AOI22_X1 U465 ( .A1(n787), .A2(\REGISTERS[18][22] ), .B1(n786), .B2(
        \REGISTERS[19][22] ), .ZN(n467) );
  AOI22_X1 U466 ( .A1(n789), .A2(\REGISTERS[20][22] ), .B1(n788), .B2(
        \REGISTERS[21][22] ), .ZN(n466) );
  AOI22_X1 U467 ( .A1(n791), .A2(\REGISTERS[4][22] ), .B1(n790), .B2(
        \REGISTERS[2][22] ), .ZN(n465) );
  AOI22_X1 U468 ( .A1(n793), .A2(\REGISTERS[26][22] ), .B1(n792), .B2(
        \REGISTERS[27][22] ), .ZN(n451) );
  AOI22_X1 U469 ( .A1(n795), .A2(\REGISTERS[28][22] ), .B1(n794), .B2(
        \REGISTERS[29][22] ), .ZN(n450) );
  AOI22_X1 U470 ( .A1(n797), .A2(\REGISTERS[30][22] ), .B1(n796), .B2(
        \REGISTERS[7][22] ), .ZN(n449) );
  AOI22_X1 U471 ( .A1(n799), .A2(\REGISTERS[5][22] ), .B1(n798), .B2(
        \REGISTERS[3][22] ), .ZN(n448) );
  NAND4_X1 U472 ( .A1(n451), .A2(n450), .A3(n449), .A4(n448), .ZN(n463) );
  AOI22_X1 U473 ( .A1(n805), .A2(\REGISTERS[9][22] ), .B1(n804), .B2(
        \REGISTERS[10][22] ), .ZN(n455) );
  AOI22_X1 U474 ( .A1(n807), .A2(\REGISTERS[11][22] ), .B1(n806), .B2(
        \REGISTERS[12][22] ), .ZN(n454) );
  AOI22_X1 U475 ( .A1(n809), .A2(\REGISTERS[13][22] ), .B1(n808), .B2(
        \REGISTERS[14][22] ), .ZN(n453) );
  AOI22_X1 U476 ( .A1(n811), .A2(\REGISTERS[15][22] ), .B1(n810), .B2(
        \REGISTERS[17][22] ), .ZN(n452) );
  NAND4_X1 U477 ( .A1(n455), .A2(n454), .A3(n453), .A4(n452), .ZN(n462) );
  AOI22_X1 U478 ( .A1(n817), .A2(\REGISTERS[31][22] ), .B1(n816), .B2(
        \REGISTERS[22][22] ), .ZN(n456) );
  OAI21_X1 U479 ( .B1(n819), .B2(n52), .A(n456), .ZN(n461) );
  AOI22_X1 U480 ( .A1(n821), .A2(\REGISTERS[24][22] ), .B1(n820), .B2(
        \REGISTERS[25][22] ), .ZN(n459) );
  AOI22_X1 U481 ( .A1(n823), .A2(\REGISTERS[8][22] ), .B1(n822), .B2(
        \REGISTERS[23][22] ), .ZN(n458) );
  AOI22_X1 U482 ( .A1(n825), .A2(\REGISTERS[16][22] ), .B1(n824), .B2(
        \REGISTERS[1][22] ), .ZN(n457) );
  NAND3_X1 U483 ( .A1(n459), .A2(n458), .A3(n457), .ZN(n460) );
  NOR4_X1 U484 ( .A1(n463), .A2(n462), .A3(n461), .A4(n460), .ZN(n464) );
  NAND4_X1 U485 ( .A1(n467), .A2(n466), .A3(n465), .A4(n464), .ZN(OUT1[22]) );
  AOI22_X1 U486 ( .A1(n71), .A2(\REGISTERS[18][23] ), .B1(n70), .B2(
        \REGISTERS[19][23] ), .ZN(n487) );
  AOI22_X1 U487 ( .A1(n73), .A2(\REGISTERS[20][23] ), .B1(n72), .B2(
        \REGISTERS[21][23] ), .ZN(n486) );
  AOI22_X1 U488 ( .A1(n791), .A2(\REGISTERS[4][23] ), .B1(n74), .B2(
        \REGISTERS[2][23] ), .ZN(n485) );
  AOI22_X1 U489 ( .A1(n77), .A2(\REGISTERS[26][23] ), .B1(n76), .B2(
        \REGISTERS[27][23] ), .ZN(n471) );
  AOI22_X1 U490 ( .A1(n79), .A2(\REGISTERS[28][23] ), .B1(n78), .B2(
        \REGISTERS[29][23] ), .ZN(n470) );
  AOI22_X1 U491 ( .A1(n81), .A2(\REGISTERS[30][23] ), .B1(n80), .B2(
        \REGISTERS[7][23] ), .ZN(n469) );
  AOI22_X1 U492 ( .A1(n83), .A2(\REGISTERS[5][23] ), .B1(n82), .B2(
        \REGISTERS[3][23] ), .ZN(n468) );
  NAND4_X1 U493 ( .A1(n471), .A2(n470), .A3(n469), .A4(n468), .ZN(n483) );
  AOI22_X1 U494 ( .A1(n85), .A2(\REGISTERS[9][23] ), .B1(n84), .B2(
        \REGISTERS[10][23] ), .ZN(n475) );
  AOI22_X1 U495 ( .A1(n87), .A2(\REGISTERS[11][23] ), .B1(n86), .B2(
        \REGISTERS[12][23] ), .ZN(n474) );
  AOI22_X1 U496 ( .A1(n89), .A2(\REGISTERS[13][23] ), .B1(n88), .B2(
        \REGISTERS[14][23] ), .ZN(n473) );
  AOI22_X1 U497 ( .A1(n91), .A2(\REGISTERS[15][23] ), .B1(n90), .B2(
        \REGISTERS[17][23] ), .ZN(n472) );
  NAND4_X1 U498 ( .A1(n475), .A2(n474), .A3(n473), .A4(n472), .ZN(n482) );
  AOI22_X1 U499 ( .A1(n93), .A2(\REGISTERS[31][23] ), .B1(n92), .B2(
        \REGISTERS[22][23] ), .ZN(n476) );
  OAI21_X1 U500 ( .B1(n819), .B2(n53), .A(n476), .ZN(n481) );
  AOI22_X1 U501 ( .A1(n95), .A2(\REGISTERS[24][23] ), .B1(n94), .B2(
        \REGISTERS[25][23] ), .ZN(n479) );
  AOI22_X1 U502 ( .A1(n97), .A2(\REGISTERS[8][23] ), .B1(n96), .B2(
        \REGISTERS[23][23] ), .ZN(n478) );
  AOI22_X1 U503 ( .A1(n825), .A2(\REGISTERS[16][23] ), .B1(n98), .B2(
        \REGISTERS[1][23] ), .ZN(n477) );
  NAND3_X1 U504 ( .A1(n479), .A2(n478), .A3(n477), .ZN(n480) );
  NOR4_X1 U505 ( .A1(n483), .A2(n482), .A3(n481), .A4(n480), .ZN(n484) );
  NAND4_X1 U506 ( .A1(n487), .A2(n486), .A3(n485), .A4(n484), .ZN(OUT1[23]) );
  AOI22_X1 U507 ( .A1(n71), .A2(\REGISTERS[18][24] ), .B1(n70), .B2(
        \REGISTERS[19][24] ), .ZN(n507) );
  AOI22_X1 U508 ( .A1(n73), .A2(\REGISTERS[20][24] ), .B1(n72), .B2(
        \REGISTERS[21][24] ), .ZN(n506) );
  AOI22_X1 U509 ( .A1(n75), .A2(\REGISTERS[4][24] ), .B1(n74), .B2(
        \REGISTERS[2][24] ), .ZN(n505) );
  AOI22_X1 U510 ( .A1(n77), .A2(\REGISTERS[26][24] ), .B1(n76), .B2(
        \REGISTERS[27][24] ), .ZN(n491) );
  AOI22_X1 U511 ( .A1(n79), .A2(\REGISTERS[28][24] ), .B1(n78), .B2(
        \REGISTERS[29][24] ), .ZN(n490) );
  AOI22_X1 U512 ( .A1(n81), .A2(\REGISTERS[30][24] ), .B1(n80), .B2(
        \REGISTERS[7][24] ), .ZN(n489) );
  AOI22_X1 U513 ( .A1(n83), .A2(\REGISTERS[5][24] ), .B1(n82), .B2(
        \REGISTERS[3][24] ), .ZN(n488) );
  NAND4_X1 U514 ( .A1(n491), .A2(n490), .A3(n489), .A4(n488), .ZN(n503) );
  AOI22_X1 U515 ( .A1(n85), .A2(\REGISTERS[9][24] ), .B1(n84), .B2(
        \REGISTERS[10][24] ), .ZN(n495) );
  AOI22_X1 U516 ( .A1(n87), .A2(\REGISTERS[11][24] ), .B1(n86), .B2(
        \REGISTERS[12][24] ), .ZN(n494) );
  AOI22_X1 U517 ( .A1(n89), .A2(\REGISTERS[13][24] ), .B1(n88), .B2(
        \REGISTERS[14][24] ), .ZN(n493) );
  AOI22_X1 U518 ( .A1(n91), .A2(\REGISTERS[15][24] ), .B1(n90), .B2(
        \REGISTERS[17][24] ), .ZN(n492) );
  NAND4_X1 U519 ( .A1(n495), .A2(n494), .A3(n493), .A4(n492), .ZN(n502) );
  AOI22_X1 U520 ( .A1(n93), .A2(\REGISTERS[31][24] ), .B1(n92), .B2(
        \REGISTERS[22][24] ), .ZN(n496) );
  OAI21_X1 U521 ( .B1(n819), .B2(n54), .A(n496), .ZN(n501) );
  AOI22_X1 U522 ( .A1(n95), .A2(\REGISTERS[24][24] ), .B1(n94), .B2(
        \REGISTERS[25][24] ), .ZN(n499) );
  AOI22_X1 U523 ( .A1(n97), .A2(\REGISTERS[8][24] ), .B1(n96), .B2(
        \REGISTERS[23][24] ), .ZN(n498) );
  AOI22_X1 U524 ( .A1(n825), .A2(\REGISTERS[16][24] ), .B1(n98), .B2(
        \REGISTERS[1][24] ), .ZN(n497) );
  NAND3_X1 U525 ( .A1(n499), .A2(n498), .A3(n497), .ZN(n500) );
  NOR4_X1 U526 ( .A1(n503), .A2(n502), .A3(n501), .A4(n500), .ZN(n504) );
  NAND4_X1 U527 ( .A1(n507), .A2(n506), .A3(n505), .A4(n504), .ZN(OUT1[24]) );
  AOI22_X1 U528 ( .A1(n71), .A2(\REGISTERS[18][25] ), .B1(n70), .B2(
        \REGISTERS[19][25] ), .ZN(n527) );
  AOI22_X1 U529 ( .A1(n73), .A2(\REGISTERS[20][25] ), .B1(n72), .B2(
        \REGISTERS[21][25] ), .ZN(n526) );
  AOI22_X1 U530 ( .A1(n75), .A2(\REGISTERS[4][25] ), .B1(n74), .B2(
        \REGISTERS[2][25] ), .ZN(n525) );
  AOI22_X1 U531 ( .A1(n793), .A2(\REGISTERS[26][25] ), .B1(n792), .B2(
        \REGISTERS[27][25] ), .ZN(n511) );
  AOI22_X1 U532 ( .A1(n795), .A2(\REGISTERS[28][25] ), .B1(n78), .B2(
        \REGISTERS[29][25] ), .ZN(n510) );
  AOI22_X1 U533 ( .A1(n797), .A2(\REGISTERS[30][25] ), .B1(n796), .B2(
        \REGISTERS[7][25] ), .ZN(n509) );
  AOI22_X1 U534 ( .A1(n799), .A2(\REGISTERS[5][25] ), .B1(n82), .B2(
        \REGISTERS[3][25] ), .ZN(n508) );
  NAND4_X1 U535 ( .A1(n511), .A2(n510), .A3(n509), .A4(n508), .ZN(n523) );
  AOI22_X1 U536 ( .A1(n805), .A2(\REGISTERS[9][25] ), .B1(n804), .B2(
        \REGISTERS[10][25] ), .ZN(n515) );
  AOI22_X1 U537 ( .A1(n807), .A2(\REGISTERS[11][25] ), .B1(n806), .B2(
        \REGISTERS[12][25] ), .ZN(n514) );
  AOI22_X1 U538 ( .A1(n809), .A2(\REGISTERS[13][25] ), .B1(n808), .B2(
        \REGISTERS[14][25] ), .ZN(n513) );
  AOI22_X1 U539 ( .A1(n811), .A2(\REGISTERS[15][25] ), .B1(n810), .B2(
        \REGISTERS[17][25] ), .ZN(n512) );
  NAND4_X1 U540 ( .A1(n515), .A2(n514), .A3(n513), .A4(n512), .ZN(n522) );
  AOI22_X1 U541 ( .A1(n817), .A2(\REGISTERS[31][25] ), .B1(n816), .B2(
        \REGISTERS[22][25] ), .ZN(n516) );
  OAI21_X1 U542 ( .B1(n819), .B2(n55), .A(n516), .ZN(n521) );
  AOI22_X1 U543 ( .A1(n821), .A2(\REGISTERS[24][25] ), .B1(n820), .B2(
        \REGISTERS[25][25] ), .ZN(n519) );
  AOI22_X1 U544 ( .A1(n97), .A2(\REGISTERS[8][25] ), .B1(n822), .B2(
        \REGISTERS[23][25] ), .ZN(n518) );
  AOI22_X1 U545 ( .A1(n825), .A2(\REGISTERS[16][25] ), .B1(n98), .B2(
        \REGISTERS[1][25] ), .ZN(n517) );
  NAND3_X1 U546 ( .A1(n519), .A2(n518), .A3(n517), .ZN(n520) );
  NOR4_X1 U547 ( .A1(n523), .A2(n522), .A3(n521), .A4(n520), .ZN(n524) );
  NAND4_X1 U548 ( .A1(n527), .A2(n526), .A3(n525), .A4(n524), .ZN(OUT1[25]) );
  AOI22_X1 U549 ( .A1(n787), .A2(\REGISTERS[18][26] ), .B1(n786), .B2(
        \REGISTERS[19][26] ), .ZN(n547) );
  AOI22_X1 U550 ( .A1(n789), .A2(\REGISTERS[20][26] ), .B1(n788), .B2(
        \REGISTERS[21][26] ), .ZN(n546) );
  AOI22_X1 U551 ( .A1(n791), .A2(\REGISTERS[4][26] ), .B1(n790), .B2(
        \REGISTERS[2][26] ), .ZN(n545) );
  AOI22_X1 U552 ( .A1(n793), .A2(\REGISTERS[26][26] ), .B1(n792), .B2(
        \REGISTERS[27][26] ), .ZN(n531) );
  AOI22_X1 U553 ( .A1(n795), .A2(\REGISTERS[28][26] ), .B1(n794), .B2(
        \REGISTERS[29][26] ), .ZN(n530) );
  AOI22_X1 U554 ( .A1(n797), .A2(\REGISTERS[30][26] ), .B1(n796), .B2(
        \REGISTERS[7][26] ), .ZN(n529) );
  AOI22_X1 U555 ( .A1(n799), .A2(\REGISTERS[5][26] ), .B1(n798), .B2(
        \REGISTERS[3][26] ), .ZN(n528) );
  NAND4_X1 U556 ( .A1(n531), .A2(n530), .A3(n529), .A4(n528), .ZN(n543) );
  AOI22_X1 U557 ( .A1(n805), .A2(\REGISTERS[9][26] ), .B1(n804), .B2(
        \REGISTERS[10][26] ), .ZN(n535) );
  AOI22_X1 U558 ( .A1(n807), .A2(\REGISTERS[11][26] ), .B1(n806), .B2(
        \REGISTERS[12][26] ), .ZN(n534) );
  AOI22_X1 U559 ( .A1(n809), .A2(\REGISTERS[13][26] ), .B1(n808), .B2(
        \REGISTERS[14][26] ), .ZN(n533) );
  AOI22_X1 U560 ( .A1(n811), .A2(\REGISTERS[15][26] ), .B1(n810), .B2(
        \REGISTERS[17][26] ), .ZN(n532) );
  NAND4_X1 U561 ( .A1(n535), .A2(n534), .A3(n533), .A4(n532), .ZN(n542) );
  AOI22_X1 U562 ( .A1(n817), .A2(\REGISTERS[31][26] ), .B1(n816), .B2(
        \REGISTERS[22][26] ), .ZN(n536) );
  OAI21_X1 U563 ( .B1(n819), .B2(n56), .A(n536), .ZN(n541) );
  AOI22_X1 U564 ( .A1(n821), .A2(\REGISTERS[24][26] ), .B1(n820), .B2(
        \REGISTERS[25][26] ), .ZN(n539) );
  AOI22_X1 U565 ( .A1(n823), .A2(\REGISTERS[8][26] ), .B1(n822), .B2(
        \REGISTERS[23][26] ), .ZN(n538) );
  AOI22_X1 U566 ( .A1(n825), .A2(\REGISTERS[16][26] ), .B1(n98), .B2(
        \REGISTERS[1][26] ), .ZN(n537) );
  NAND3_X1 U567 ( .A1(n539), .A2(n538), .A3(n537), .ZN(n540) );
  NOR4_X1 U568 ( .A1(n543), .A2(n542), .A3(n541), .A4(n540), .ZN(n544) );
  NAND4_X1 U569 ( .A1(n547), .A2(n546), .A3(n545), .A4(n544), .ZN(OUT1[26]) );
  AOI22_X1 U570 ( .A1(n71), .A2(\REGISTERS[18][27] ), .B1(n70), .B2(
        \REGISTERS[19][27] ), .ZN(n567) );
  AOI22_X1 U571 ( .A1(n789), .A2(\REGISTERS[20][27] ), .B1(n72), .B2(
        \REGISTERS[21][27] ), .ZN(n566) );
  AOI22_X1 U572 ( .A1(n791), .A2(\REGISTERS[4][27] ), .B1(n790), .B2(
        \REGISTERS[2][27] ), .ZN(n565) );
  AOI22_X1 U573 ( .A1(n77), .A2(\REGISTERS[26][27] ), .B1(n76), .B2(
        \REGISTERS[27][27] ), .ZN(n551) );
  AOI22_X1 U574 ( .A1(n79), .A2(\REGISTERS[28][27] ), .B1(n78), .B2(
        \REGISTERS[29][27] ), .ZN(n550) );
  AOI22_X1 U575 ( .A1(n81), .A2(\REGISTERS[30][27] ), .B1(n80), .B2(
        \REGISTERS[7][27] ), .ZN(n549) );
  AOI22_X1 U576 ( .A1(n83), .A2(\REGISTERS[5][27] ), .B1(n798), .B2(
        \REGISTERS[3][27] ), .ZN(n548) );
  NAND4_X1 U577 ( .A1(n551), .A2(n550), .A3(n549), .A4(n548), .ZN(n563) );
  AOI22_X1 U578 ( .A1(n805), .A2(\REGISTERS[9][27] ), .B1(n804), .B2(
        \REGISTERS[10][27] ), .ZN(n555) );
  AOI22_X1 U579 ( .A1(n87), .A2(\REGISTERS[11][27] ), .B1(n806), .B2(
        \REGISTERS[12][27] ), .ZN(n554) );
  AOI22_X1 U580 ( .A1(n89), .A2(\REGISTERS[13][27] ), .B1(n808), .B2(
        \REGISTERS[14][27] ), .ZN(n553) );
  AOI22_X1 U581 ( .A1(n811), .A2(\REGISTERS[15][27] ), .B1(n90), .B2(
        \REGISTERS[17][27] ), .ZN(n552) );
  NAND4_X1 U582 ( .A1(n555), .A2(n554), .A3(n553), .A4(n552), .ZN(n562) );
  AOI22_X1 U583 ( .A1(n93), .A2(\REGISTERS[31][27] ), .B1(n92), .B2(
        \REGISTERS[22][27] ), .ZN(n556) );
  OAI21_X1 U584 ( .B1(n819), .B2(n57), .A(n556), .ZN(n561) );
  AOI22_X1 U585 ( .A1(n95), .A2(\REGISTERS[24][27] ), .B1(n94), .B2(
        \REGISTERS[25][27] ), .ZN(n559) );
  AOI22_X1 U586 ( .A1(n97), .A2(\REGISTERS[8][27] ), .B1(n96), .B2(
        \REGISTERS[23][27] ), .ZN(n558) );
  AOI22_X1 U587 ( .A1(n825), .A2(\REGISTERS[16][27] ), .B1(n98), .B2(
        \REGISTERS[1][27] ), .ZN(n557) );
  NAND3_X1 U588 ( .A1(n559), .A2(n558), .A3(n557), .ZN(n560) );
  NOR4_X1 U589 ( .A1(n563), .A2(n562), .A3(n561), .A4(n560), .ZN(n564) );
  NAND4_X1 U590 ( .A1(n567), .A2(n566), .A3(n565), .A4(n564), .ZN(OUT1[27]) );
  AOI22_X1 U591 ( .A1(n71), .A2(\REGISTERS[18][28] ), .B1(n70), .B2(
        \REGISTERS[19][28] ), .ZN(n587) );
  AOI22_X1 U592 ( .A1(n73), .A2(\REGISTERS[20][28] ), .B1(n72), .B2(
        \REGISTERS[21][28] ), .ZN(n586) );
  AOI22_X1 U593 ( .A1(n75), .A2(\REGISTERS[4][28] ), .B1(n74), .B2(
        \REGISTERS[2][28] ), .ZN(n585) );
  AOI22_X1 U594 ( .A1(n77), .A2(\REGISTERS[26][28] ), .B1(n76), .B2(
        \REGISTERS[27][28] ), .ZN(n571) );
  AOI22_X1 U595 ( .A1(n79), .A2(\REGISTERS[28][28] ), .B1(n78), .B2(
        \REGISTERS[29][28] ), .ZN(n570) );
  AOI22_X1 U596 ( .A1(n81), .A2(\REGISTERS[30][28] ), .B1(n80), .B2(
        \REGISTERS[7][28] ), .ZN(n569) );
  AOI22_X1 U597 ( .A1(n83), .A2(\REGISTERS[5][28] ), .B1(n82), .B2(
        \REGISTERS[3][28] ), .ZN(n568) );
  NAND4_X1 U598 ( .A1(n571), .A2(n570), .A3(n569), .A4(n568), .ZN(n583) );
  AOI22_X1 U599 ( .A1(n85), .A2(\REGISTERS[9][28] ), .B1(n84), .B2(
        \REGISTERS[10][28] ), .ZN(n575) );
  AOI22_X1 U600 ( .A1(n87), .A2(\REGISTERS[11][28] ), .B1(n86), .B2(
        \REGISTERS[12][28] ), .ZN(n574) );
  AOI22_X1 U601 ( .A1(n89), .A2(\REGISTERS[13][28] ), .B1(n88), .B2(
        \REGISTERS[14][28] ), .ZN(n573) );
  AOI22_X1 U602 ( .A1(n91), .A2(\REGISTERS[15][28] ), .B1(n90), .B2(
        \REGISTERS[17][28] ), .ZN(n572) );
  NAND4_X1 U603 ( .A1(n575), .A2(n574), .A3(n573), .A4(n572), .ZN(n582) );
  AOI22_X1 U604 ( .A1(n93), .A2(\REGISTERS[31][28] ), .B1(n92), .B2(
        \REGISTERS[22][28] ), .ZN(n576) );
  OAI21_X1 U605 ( .B1(n819), .B2(n58), .A(n576), .ZN(n581) );
  AOI22_X1 U606 ( .A1(n95), .A2(\REGISTERS[24][28] ), .B1(n94), .B2(
        \REGISTERS[25][28] ), .ZN(n579) );
  AOI22_X1 U607 ( .A1(n97), .A2(\REGISTERS[8][28] ), .B1(n96), .B2(
        \REGISTERS[23][28] ), .ZN(n578) );
  AOI22_X1 U608 ( .A1(n825), .A2(\REGISTERS[16][28] ), .B1(n98), .B2(
        \REGISTERS[1][28] ), .ZN(n577) );
  NAND3_X1 U609 ( .A1(n579), .A2(n578), .A3(n577), .ZN(n580) );
  NOR4_X1 U610 ( .A1(n583), .A2(n582), .A3(n581), .A4(n580), .ZN(n584) );
  NAND4_X1 U611 ( .A1(n587), .A2(n586), .A3(n585), .A4(n584), .ZN(OUT1[28]) );
  AOI22_X1 U612 ( .A1(n71), .A2(\REGISTERS[18][29] ), .B1(n70), .B2(
        \REGISTERS[19][29] ), .ZN(n607) );
  AOI22_X1 U613 ( .A1(n73), .A2(\REGISTERS[20][29] ), .B1(n72), .B2(
        \REGISTERS[21][29] ), .ZN(n606) );
  AOI22_X1 U614 ( .A1(n75), .A2(\REGISTERS[4][29] ), .B1(n74), .B2(
        \REGISTERS[2][29] ), .ZN(n605) );
  AOI22_X1 U615 ( .A1(n77), .A2(\REGISTERS[26][29] ), .B1(n76), .B2(
        \REGISTERS[27][29] ), .ZN(n591) );
  AOI22_X1 U616 ( .A1(n79), .A2(\REGISTERS[28][29] ), .B1(n78), .B2(
        \REGISTERS[29][29] ), .ZN(n590) );
  AOI22_X1 U617 ( .A1(n797), .A2(\REGISTERS[30][29] ), .B1(n796), .B2(
        \REGISTERS[7][29] ), .ZN(n589) );
  AOI22_X1 U618 ( .A1(n799), .A2(\REGISTERS[5][29] ), .B1(n82), .B2(
        \REGISTERS[3][29] ), .ZN(n588) );
  NAND4_X1 U619 ( .A1(n591), .A2(n590), .A3(n589), .A4(n588), .ZN(n603) );
  AOI22_X1 U620 ( .A1(n85), .A2(\REGISTERS[9][29] ), .B1(n84), .B2(
        \REGISTERS[10][29] ), .ZN(n595) );
  AOI22_X1 U621 ( .A1(n87), .A2(\REGISTERS[11][29] ), .B1(n86), .B2(
        \REGISTERS[12][29] ), .ZN(n594) );
  AOI22_X1 U622 ( .A1(n89), .A2(\REGISTERS[13][29] ), .B1(n88), .B2(
        \REGISTERS[14][29] ), .ZN(n593) );
  AOI22_X1 U623 ( .A1(n91), .A2(\REGISTERS[15][29] ), .B1(n810), .B2(
        \REGISTERS[17][29] ), .ZN(n592) );
  NAND4_X1 U624 ( .A1(n595), .A2(n594), .A3(n593), .A4(n592), .ZN(n602) );
  AOI22_X1 U625 ( .A1(n817), .A2(\REGISTERS[31][29] ), .B1(n816), .B2(
        \REGISTERS[22][29] ), .ZN(n596) );
  OAI21_X1 U626 ( .B1(n819), .B2(n59), .A(n596), .ZN(n601) );
  AOI22_X1 U627 ( .A1(n95), .A2(\REGISTERS[24][29] ), .B1(n820), .B2(
        \REGISTERS[25][29] ), .ZN(n599) );
  AOI22_X1 U628 ( .A1(n97), .A2(\REGISTERS[8][29] ), .B1(n822), .B2(
        \REGISTERS[23][29] ), .ZN(n598) );
  AOI22_X1 U629 ( .A1(n825), .A2(\REGISTERS[16][29] ), .B1(n98), .B2(
        \REGISTERS[1][29] ), .ZN(n597) );
  NAND3_X1 U630 ( .A1(n599), .A2(n598), .A3(n597), .ZN(n600) );
  NOR4_X1 U631 ( .A1(n603), .A2(n602), .A3(n601), .A4(n600), .ZN(n604) );
  NAND4_X1 U632 ( .A1(n607), .A2(n606), .A3(n605), .A4(n604), .ZN(OUT1[29]) );
  AOI22_X1 U633 ( .A1(n71), .A2(\REGISTERS[18][2] ), .B1(n70), .B2(
        \REGISTERS[19][2] ), .ZN(n627) );
  AOI22_X1 U634 ( .A1(n73), .A2(\REGISTERS[20][2] ), .B1(n72), .B2(
        \REGISTERS[21][2] ), .ZN(n626) );
  AOI22_X1 U635 ( .A1(n75), .A2(\REGISTERS[4][2] ), .B1(n74), .B2(
        \REGISTERS[2][2] ), .ZN(n625) );
  AOI22_X1 U636 ( .A1(n77), .A2(\REGISTERS[26][2] ), .B1(n76), .B2(
        \REGISTERS[27][2] ), .ZN(n611) );
  AOI22_X1 U637 ( .A1(n79), .A2(\REGISTERS[28][2] ), .B1(n78), .B2(
        \REGISTERS[29][2] ), .ZN(n610) );
  AOI22_X1 U638 ( .A1(n81), .A2(\REGISTERS[30][2] ), .B1(n80), .B2(
        \REGISTERS[7][2] ), .ZN(n609) );
  AOI22_X1 U639 ( .A1(n83), .A2(\REGISTERS[5][2] ), .B1(n82), .B2(
        \REGISTERS[3][2] ), .ZN(n608) );
  NAND4_X1 U640 ( .A1(n611), .A2(n610), .A3(n609), .A4(n608), .ZN(n623) );
  AOI22_X1 U641 ( .A1(n85), .A2(\REGISTERS[9][2] ), .B1(n84), .B2(
        \REGISTERS[10][2] ), .ZN(n615) );
  AOI22_X1 U642 ( .A1(n87), .A2(\REGISTERS[11][2] ), .B1(n86), .B2(
        \REGISTERS[12][2] ), .ZN(n614) );
  AOI22_X1 U643 ( .A1(n89), .A2(\REGISTERS[13][2] ), .B1(n88), .B2(
        \REGISTERS[14][2] ), .ZN(n613) );
  AOI22_X1 U644 ( .A1(n91), .A2(\REGISTERS[15][2] ), .B1(n90), .B2(
        \REGISTERS[17][2] ), .ZN(n612) );
  NAND4_X1 U645 ( .A1(n615), .A2(n614), .A3(n613), .A4(n612), .ZN(n622) );
  AOI22_X1 U646 ( .A1(n93), .A2(\REGISTERS[31][2] ), .B1(n92), .B2(
        \REGISTERS[22][2] ), .ZN(n616) );
  OAI21_X1 U647 ( .B1(n819), .B2(n60), .A(n616), .ZN(n621) );
  AOI22_X1 U648 ( .A1(n95), .A2(\REGISTERS[24][2] ), .B1(n94), .B2(
        \REGISTERS[25][2] ), .ZN(n619) );
  AOI22_X1 U649 ( .A1(n97), .A2(\REGISTERS[8][2] ), .B1(n96), .B2(
        \REGISTERS[23][2] ), .ZN(n618) );
  AOI22_X1 U650 ( .A1(n825), .A2(\REGISTERS[16][2] ), .B1(n98), .B2(
        \REGISTERS[1][2] ), .ZN(n617) );
  NAND3_X1 U651 ( .A1(n619), .A2(n618), .A3(n617), .ZN(n620) );
  NOR4_X1 U652 ( .A1(n623), .A2(n622), .A3(n621), .A4(n620), .ZN(n624) );
  NAND4_X1 U653 ( .A1(n627), .A2(n626), .A3(n625), .A4(n624), .ZN(OUT1[2]) );
  AOI22_X1 U654 ( .A1(n75), .A2(\REGISTERS[4][30] ), .B1(n74), .B2(
        \REGISTERS[2][30] ), .ZN(n645) );
  AOI22_X1 U655 ( .A1(n77), .A2(\REGISTERS[26][30] ), .B1(n76), .B2(
        \REGISTERS[27][30] ), .ZN(n631) );
  AOI22_X1 U656 ( .A1(n79), .A2(\REGISTERS[28][30] ), .B1(n78), .B2(
        \REGISTERS[29][30] ), .ZN(n630) );
  AOI22_X1 U657 ( .A1(n81), .A2(\REGISTERS[30][30] ), .B1(n80), .B2(
        \REGISTERS[7][30] ), .ZN(n629) );
  AOI22_X1 U658 ( .A1(n83), .A2(\REGISTERS[5][30] ), .B1(n82), .B2(
        \REGISTERS[3][30] ), .ZN(n628) );
  NAND4_X1 U659 ( .A1(n631), .A2(n630), .A3(n629), .A4(n628), .ZN(n643) );
  AOI22_X1 U660 ( .A1(n85), .A2(\REGISTERS[9][30] ), .B1(n84), .B2(
        \REGISTERS[10][30] ), .ZN(n635) );
  AOI22_X1 U661 ( .A1(n87), .A2(\REGISTERS[11][30] ), .B1(n86), .B2(
        \REGISTERS[12][30] ), .ZN(n634) );
  AOI22_X1 U662 ( .A1(n89), .A2(\REGISTERS[13][30] ), .B1(n88), .B2(
        \REGISTERS[14][30] ), .ZN(n633) );
  AOI22_X1 U663 ( .A1(n91), .A2(\REGISTERS[15][30] ), .B1(n90), .B2(
        \REGISTERS[17][30] ), .ZN(n632) );
  NAND4_X1 U664 ( .A1(n635), .A2(n634), .A3(n633), .A4(n632), .ZN(n642) );
  AOI22_X1 U665 ( .A1(n93), .A2(\REGISTERS[31][30] ), .B1(n92), .B2(
        \REGISTERS[22][30] ), .ZN(n636) );
  OAI21_X1 U666 ( .B1(n819), .B2(n61), .A(n636), .ZN(n641) );
  AOI22_X1 U667 ( .A1(n95), .A2(\REGISTERS[24][30] ), .B1(n94), .B2(
        \REGISTERS[25][30] ), .ZN(n639) );
  AOI22_X1 U668 ( .A1(n97), .A2(\REGISTERS[8][30] ), .B1(n96), .B2(
        \REGISTERS[23][30] ), .ZN(n638) );
  AOI22_X1 U669 ( .A1(n825), .A2(\REGISTERS[16][30] ), .B1(n98), .B2(
        \REGISTERS[1][30] ), .ZN(n637) );
  NAND3_X1 U670 ( .A1(n639), .A2(n638), .A3(n637), .ZN(n640) );
  NOR4_X1 U671 ( .A1(n643), .A2(n642), .A3(n641), .A4(n640), .ZN(n644) );
  AOI22_X1 U672 ( .A1(n71), .A2(\REGISTERS[18][31] ), .B1(n70), .B2(
        \REGISTERS[19][31] ), .ZN(n665) );
  AOI22_X1 U673 ( .A1(n73), .A2(\REGISTERS[20][31] ), .B1(n72), .B2(
        \REGISTERS[21][31] ), .ZN(n664) );
  AOI22_X1 U674 ( .A1(n75), .A2(\REGISTERS[4][31] ), .B1(n74), .B2(
        \REGISTERS[2][31] ), .ZN(n663) );
  AOI22_X1 U675 ( .A1(n77), .A2(\REGISTERS[26][31] ), .B1(n76), .B2(
        \REGISTERS[27][31] ), .ZN(n649) );
  AOI22_X1 U676 ( .A1(n79), .A2(\REGISTERS[28][31] ), .B1(n78), .B2(
        \REGISTERS[29][31] ), .ZN(n648) );
  AOI22_X1 U677 ( .A1(n81), .A2(\REGISTERS[30][31] ), .B1(n80), .B2(
        \REGISTERS[7][31] ), .ZN(n647) );
  AOI22_X1 U678 ( .A1(n83), .A2(\REGISTERS[5][31] ), .B1(n82), .B2(
        \REGISTERS[3][31] ), .ZN(n646) );
  NAND4_X1 U679 ( .A1(n649), .A2(n648), .A3(n647), .A4(n646), .ZN(n661) );
  AOI22_X1 U680 ( .A1(n85), .A2(\REGISTERS[9][31] ), .B1(n84), .B2(
        \REGISTERS[10][31] ), .ZN(n653) );
  AOI22_X1 U681 ( .A1(n87), .A2(\REGISTERS[11][31] ), .B1(n86), .B2(
        \REGISTERS[12][31] ), .ZN(n652) );
  AOI22_X1 U682 ( .A1(n89), .A2(\REGISTERS[13][31] ), .B1(n88), .B2(
        \REGISTERS[14][31] ), .ZN(n651) );
  AOI22_X1 U683 ( .A1(n91), .A2(\REGISTERS[15][31] ), .B1(n90), .B2(
        \REGISTERS[17][31] ), .ZN(n650) );
  NAND4_X1 U684 ( .A1(n653), .A2(n652), .A3(n651), .A4(n650), .ZN(n660) );
  AOI22_X1 U685 ( .A1(n93), .A2(\REGISTERS[31][31] ), .B1(n92), .B2(
        \REGISTERS[22][31] ), .ZN(n654) );
  OAI21_X1 U686 ( .B1(n819), .B2(n62), .A(n654), .ZN(n659) );
  AOI22_X1 U687 ( .A1(n95), .A2(\REGISTERS[24][31] ), .B1(n94), .B2(
        \REGISTERS[25][31] ), .ZN(n657) );
  AOI22_X1 U688 ( .A1(n97), .A2(\REGISTERS[8][31] ), .B1(n96), .B2(
        \REGISTERS[23][31] ), .ZN(n656) );
  AOI22_X1 U689 ( .A1(n825), .A2(\REGISTERS[16][31] ), .B1(n98), .B2(
        \REGISTERS[1][31] ), .ZN(n655) );
  NAND3_X1 U690 ( .A1(n657), .A2(n656), .A3(n655), .ZN(n658) );
  NOR4_X1 U691 ( .A1(n661), .A2(n660), .A3(n659), .A4(n658), .ZN(n662) );
  NAND4_X1 U692 ( .A1(n665), .A2(n664), .A3(n663), .A4(n662), .ZN(OUT1[31]) );
  AOI22_X1 U693 ( .A1(n71), .A2(\REGISTERS[18][3] ), .B1(n70), .B2(
        \REGISTERS[19][3] ), .ZN(n685) );
  AOI22_X1 U694 ( .A1(n73), .A2(\REGISTERS[20][3] ), .B1(n72), .B2(
        \REGISTERS[21][3] ), .ZN(n684) );
  AOI22_X1 U695 ( .A1(n75), .A2(\REGISTERS[4][3] ), .B1(n74), .B2(
        \REGISTERS[2][3] ), .ZN(n683) );
  AOI22_X1 U696 ( .A1(n77), .A2(\REGISTERS[26][3] ), .B1(n76), .B2(
        \REGISTERS[27][3] ), .ZN(n669) );
  AOI22_X1 U697 ( .A1(n79), .A2(\REGISTERS[28][3] ), .B1(n78), .B2(
        \REGISTERS[29][3] ), .ZN(n668) );
  AOI22_X1 U698 ( .A1(n81), .A2(\REGISTERS[30][3] ), .B1(n80), .B2(
        \REGISTERS[7][3] ), .ZN(n667) );
  AOI22_X1 U699 ( .A1(n83), .A2(\REGISTERS[5][3] ), .B1(n82), .B2(
        \REGISTERS[3][3] ), .ZN(n666) );
  NAND4_X1 U700 ( .A1(n669), .A2(n668), .A3(n667), .A4(n666), .ZN(n681) );
  AOI22_X1 U701 ( .A1(n85), .A2(\REGISTERS[9][3] ), .B1(n84), .B2(
        \REGISTERS[10][3] ), .ZN(n673) );
  AOI22_X1 U702 ( .A1(n87), .A2(\REGISTERS[11][3] ), .B1(n86), .B2(
        \REGISTERS[12][3] ), .ZN(n672) );
  AOI22_X1 U703 ( .A1(n89), .A2(\REGISTERS[13][3] ), .B1(n88), .B2(
        \REGISTERS[14][3] ), .ZN(n671) );
  AOI22_X1 U704 ( .A1(n91), .A2(\REGISTERS[15][3] ), .B1(n90), .B2(
        \REGISTERS[17][3] ), .ZN(n670) );
  NAND4_X1 U705 ( .A1(n673), .A2(n672), .A3(n671), .A4(n670), .ZN(n680) );
  AOI22_X1 U706 ( .A1(n93), .A2(\REGISTERS[31][3] ), .B1(n92), .B2(
        \REGISTERS[22][3] ), .ZN(n674) );
  OAI21_X1 U707 ( .B1(n819), .B2(n63), .A(n674), .ZN(n679) );
  AOI22_X1 U708 ( .A1(n95), .A2(\REGISTERS[24][3] ), .B1(n94), .B2(
        \REGISTERS[25][3] ), .ZN(n677) );
  AOI22_X1 U709 ( .A1(n97), .A2(\REGISTERS[8][3] ), .B1(n96), .B2(
        \REGISTERS[23][3] ), .ZN(n676) );
  AOI22_X1 U710 ( .A1(n825), .A2(\REGISTERS[16][3] ), .B1(n98), .B2(
        \REGISTERS[1][3] ), .ZN(n675) );
  NAND3_X1 U711 ( .A1(n677), .A2(n676), .A3(n675), .ZN(n678) );
  NOR4_X1 U712 ( .A1(n681), .A2(n680), .A3(n679), .A4(n678), .ZN(n682) );
  NAND4_X1 U713 ( .A1(n685), .A2(n684), .A3(n683), .A4(n682), .ZN(OUT1[3]) );
  AOI22_X1 U714 ( .A1(n71), .A2(\REGISTERS[18][4] ), .B1(n70), .B2(
        \REGISTERS[19][4] ), .ZN(n705) );
  AOI22_X1 U715 ( .A1(n73), .A2(\REGISTERS[20][4] ), .B1(n72), .B2(
        \REGISTERS[21][4] ), .ZN(n704) );
  AOI22_X1 U716 ( .A1(n75), .A2(\REGISTERS[4][4] ), .B1(n74), .B2(
        \REGISTERS[2][4] ), .ZN(n703) );
  AOI22_X1 U717 ( .A1(n77), .A2(\REGISTERS[26][4] ), .B1(n76), .B2(
        \REGISTERS[27][4] ), .ZN(n689) );
  AOI22_X1 U718 ( .A1(n79), .A2(\REGISTERS[28][4] ), .B1(n78), .B2(
        \REGISTERS[29][4] ), .ZN(n688) );
  AOI22_X1 U719 ( .A1(n81), .A2(\REGISTERS[30][4] ), .B1(n80), .B2(
        \REGISTERS[7][4] ), .ZN(n687) );
  AOI22_X1 U720 ( .A1(n83), .A2(\REGISTERS[5][4] ), .B1(n82), .B2(
        \REGISTERS[3][4] ), .ZN(n686) );
  NAND4_X1 U721 ( .A1(n689), .A2(n688), .A3(n687), .A4(n686), .ZN(n701) );
  AOI22_X1 U722 ( .A1(n85), .A2(\REGISTERS[9][4] ), .B1(n84), .B2(
        \REGISTERS[10][4] ), .ZN(n693) );
  AOI22_X1 U723 ( .A1(n87), .A2(\REGISTERS[11][4] ), .B1(n86), .B2(
        \REGISTERS[12][4] ), .ZN(n692) );
  AOI22_X1 U724 ( .A1(n89), .A2(\REGISTERS[13][4] ), .B1(n88), .B2(
        \REGISTERS[14][4] ), .ZN(n691) );
  AOI22_X1 U725 ( .A1(n91), .A2(\REGISTERS[15][4] ), .B1(n90), .B2(
        \REGISTERS[17][4] ), .ZN(n690) );
  NAND4_X1 U726 ( .A1(n693), .A2(n692), .A3(n691), .A4(n690), .ZN(n700) );
  AOI22_X1 U727 ( .A1(n93), .A2(\REGISTERS[31][4] ), .B1(n92), .B2(
        \REGISTERS[22][4] ), .ZN(n694) );
  OAI21_X1 U728 ( .B1(n819), .B2(n64), .A(n694), .ZN(n699) );
  AOI22_X1 U729 ( .A1(n95), .A2(\REGISTERS[24][4] ), .B1(n94), .B2(
        \REGISTERS[25][4] ), .ZN(n697) );
  AOI22_X1 U730 ( .A1(n97), .A2(\REGISTERS[8][4] ), .B1(n96), .B2(
        \REGISTERS[23][4] ), .ZN(n696) );
  AOI22_X1 U731 ( .A1(n825), .A2(\REGISTERS[16][4] ), .B1(n98), .B2(
        \REGISTERS[1][4] ), .ZN(n695) );
  NAND3_X1 U732 ( .A1(n697), .A2(n696), .A3(n695), .ZN(n698) );
  NOR4_X1 U733 ( .A1(n701), .A2(n700), .A3(n699), .A4(n698), .ZN(n702) );
  NAND4_X1 U734 ( .A1(n705), .A2(n704), .A3(n703), .A4(n702), .ZN(OUT1[4]) );
  AOI22_X1 U735 ( .A1(n71), .A2(\REGISTERS[18][5] ), .B1(n70), .B2(
        \REGISTERS[19][5] ), .ZN(n725) );
  AOI22_X1 U736 ( .A1(n73), .A2(\REGISTERS[20][5] ), .B1(n72), .B2(
        \REGISTERS[21][5] ), .ZN(n724) );
  AOI22_X1 U737 ( .A1(n75), .A2(\REGISTERS[4][5] ), .B1(n74), .B2(
        \REGISTERS[2][5] ), .ZN(n723) );
  AOI22_X1 U738 ( .A1(n77), .A2(\REGISTERS[26][5] ), .B1(n76), .B2(
        \REGISTERS[27][5] ), .ZN(n709) );
  AOI22_X1 U739 ( .A1(n79), .A2(\REGISTERS[28][5] ), .B1(n78), .B2(
        \REGISTERS[29][5] ), .ZN(n708) );
  AOI22_X1 U740 ( .A1(n81), .A2(\REGISTERS[30][5] ), .B1(n80), .B2(
        \REGISTERS[7][5] ), .ZN(n707) );
  AOI22_X1 U741 ( .A1(n83), .A2(\REGISTERS[5][5] ), .B1(n82), .B2(
        \REGISTERS[3][5] ), .ZN(n706) );
  NAND4_X1 U742 ( .A1(n709), .A2(n708), .A3(n707), .A4(n706), .ZN(n721) );
  AOI22_X1 U743 ( .A1(n85), .A2(\REGISTERS[9][5] ), .B1(n84), .B2(
        \REGISTERS[10][5] ), .ZN(n713) );
  AOI22_X1 U744 ( .A1(n87), .A2(\REGISTERS[11][5] ), .B1(n86), .B2(
        \REGISTERS[12][5] ), .ZN(n712) );
  AOI22_X1 U745 ( .A1(n89), .A2(\REGISTERS[13][5] ), .B1(n88), .B2(
        \REGISTERS[14][5] ), .ZN(n711) );
  AOI22_X1 U746 ( .A1(n91), .A2(\REGISTERS[15][5] ), .B1(n90), .B2(
        \REGISTERS[17][5] ), .ZN(n710) );
  NAND4_X1 U747 ( .A1(n713), .A2(n712), .A3(n711), .A4(n710), .ZN(n720) );
  AOI22_X1 U748 ( .A1(n93), .A2(\REGISTERS[31][5] ), .B1(n92), .B2(
        \REGISTERS[22][5] ), .ZN(n714) );
  OAI21_X1 U749 ( .B1(n819), .B2(n65), .A(n714), .ZN(n719) );
  AOI22_X1 U750 ( .A1(n95), .A2(\REGISTERS[24][5] ), .B1(n94), .B2(
        \REGISTERS[25][5] ), .ZN(n717) );
  AOI22_X1 U751 ( .A1(n97), .A2(\REGISTERS[8][5] ), .B1(n96), .B2(
        \REGISTERS[23][5] ), .ZN(n716) );
  AOI22_X1 U752 ( .A1(n825), .A2(\REGISTERS[16][5] ), .B1(n98), .B2(
        \REGISTERS[1][5] ), .ZN(n715) );
  NAND3_X1 U753 ( .A1(n717), .A2(n716), .A3(n715), .ZN(n718) );
  NOR4_X1 U754 ( .A1(n721), .A2(n720), .A3(n719), .A4(n718), .ZN(n722) );
  NAND4_X1 U755 ( .A1(n725), .A2(n724), .A3(n723), .A4(n722), .ZN(OUT1[5]) );
  AOI22_X1 U756 ( .A1(n71), .A2(\REGISTERS[18][6] ), .B1(n70), .B2(
        \REGISTERS[19][6] ), .ZN(n745) );
  AOI22_X1 U757 ( .A1(n73), .A2(\REGISTERS[20][6] ), .B1(n72), .B2(
        \REGISTERS[21][6] ), .ZN(n744) );
  AOI22_X1 U758 ( .A1(n75), .A2(\REGISTERS[4][6] ), .B1(n74), .B2(
        \REGISTERS[2][6] ), .ZN(n743) );
  AOI22_X1 U759 ( .A1(n77), .A2(\REGISTERS[26][6] ), .B1(n76), .B2(
        \REGISTERS[27][6] ), .ZN(n729) );
  AOI22_X1 U760 ( .A1(n79), .A2(\REGISTERS[28][6] ), .B1(n78), .B2(
        \REGISTERS[29][6] ), .ZN(n728) );
  AOI22_X1 U761 ( .A1(n81), .A2(\REGISTERS[30][6] ), .B1(n80), .B2(
        \REGISTERS[7][6] ), .ZN(n727) );
  AOI22_X1 U762 ( .A1(n83), .A2(\REGISTERS[5][6] ), .B1(n82), .B2(
        \REGISTERS[3][6] ), .ZN(n726) );
  NAND4_X1 U763 ( .A1(n729), .A2(n728), .A3(n727), .A4(n726), .ZN(n741) );
  AOI22_X1 U764 ( .A1(n85), .A2(\REGISTERS[9][6] ), .B1(n84), .B2(
        \REGISTERS[10][6] ), .ZN(n733) );
  AOI22_X1 U765 ( .A1(n87), .A2(\REGISTERS[11][6] ), .B1(n86), .B2(
        \REGISTERS[12][6] ), .ZN(n732) );
  AOI22_X1 U766 ( .A1(n89), .A2(\REGISTERS[13][6] ), .B1(n88), .B2(
        \REGISTERS[14][6] ), .ZN(n731) );
  AOI22_X1 U767 ( .A1(n91), .A2(\REGISTERS[15][6] ), .B1(n90), .B2(
        \REGISTERS[17][6] ), .ZN(n730) );
  NAND4_X1 U768 ( .A1(n733), .A2(n732), .A3(n731), .A4(n730), .ZN(n740) );
  AOI22_X1 U769 ( .A1(n93), .A2(\REGISTERS[31][6] ), .B1(n92), .B2(
        \REGISTERS[22][6] ), .ZN(n734) );
  OAI21_X1 U770 ( .B1(n819), .B2(n66), .A(n734), .ZN(n739) );
  AOI22_X1 U771 ( .A1(n95), .A2(\REGISTERS[24][6] ), .B1(n94), .B2(
        \REGISTERS[25][6] ), .ZN(n737) );
  AOI22_X1 U772 ( .A1(n97), .A2(\REGISTERS[8][6] ), .B1(n96), .B2(
        \REGISTERS[23][6] ), .ZN(n736) );
  AOI22_X1 U773 ( .A1(n825), .A2(\REGISTERS[16][6] ), .B1(n98), .B2(
        \REGISTERS[1][6] ), .ZN(n735) );
  NAND3_X1 U774 ( .A1(n737), .A2(n736), .A3(n735), .ZN(n738) );
  NOR4_X1 U775 ( .A1(n741), .A2(n740), .A3(n739), .A4(n738), .ZN(n742) );
  NAND4_X1 U776 ( .A1(n745), .A2(n744), .A3(n743), .A4(n742), .ZN(OUT1[6]) );
  AOI22_X1 U777 ( .A1(n71), .A2(\REGISTERS[18][7] ), .B1(n70), .B2(
        \REGISTERS[19][7] ), .ZN(n765) );
  AOI22_X1 U778 ( .A1(n73), .A2(\REGISTERS[20][7] ), .B1(n72), .B2(
        \REGISTERS[21][7] ), .ZN(n764) );
  AOI22_X1 U779 ( .A1(n75), .A2(\REGISTERS[4][7] ), .B1(n74), .B2(
        \REGISTERS[2][7] ), .ZN(n763) );
  AOI22_X1 U780 ( .A1(n77), .A2(\REGISTERS[26][7] ), .B1(n76), .B2(
        \REGISTERS[27][7] ), .ZN(n749) );
  AOI22_X1 U781 ( .A1(n79), .A2(\REGISTERS[28][7] ), .B1(n78), .B2(
        \REGISTERS[29][7] ), .ZN(n748) );
  AOI22_X1 U782 ( .A1(n81), .A2(\REGISTERS[30][7] ), .B1(n80), .B2(
        \REGISTERS[7][7] ), .ZN(n747) );
  AOI22_X1 U783 ( .A1(n83), .A2(\REGISTERS[5][7] ), .B1(n82), .B2(
        \REGISTERS[3][7] ), .ZN(n746) );
  NAND4_X1 U784 ( .A1(n749), .A2(n748), .A3(n747), .A4(n746), .ZN(n761) );
  AOI22_X1 U785 ( .A1(n85), .A2(\REGISTERS[9][7] ), .B1(n84), .B2(
        \REGISTERS[10][7] ), .ZN(n753) );
  AOI22_X1 U786 ( .A1(n87), .A2(\REGISTERS[11][7] ), .B1(n86), .B2(
        \REGISTERS[12][7] ), .ZN(n752) );
  AOI22_X1 U787 ( .A1(n89), .A2(\REGISTERS[13][7] ), .B1(n88), .B2(
        \REGISTERS[14][7] ), .ZN(n751) );
  AOI22_X1 U788 ( .A1(n91), .A2(\REGISTERS[15][7] ), .B1(n90), .B2(
        \REGISTERS[17][7] ), .ZN(n750) );
  NAND4_X1 U789 ( .A1(n753), .A2(n752), .A3(n751), .A4(n750), .ZN(n760) );
  AOI22_X1 U790 ( .A1(n93), .A2(\REGISTERS[31][7] ), .B1(n92), .B2(
        \REGISTERS[22][7] ), .ZN(n754) );
  OAI21_X1 U791 ( .B1(n819), .B2(n67), .A(n754), .ZN(n759) );
  AOI22_X1 U792 ( .A1(n95), .A2(\REGISTERS[24][7] ), .B1(n94), .B2(
        \REGISTERS[25][7] ), .ZN(n757) );
  AOI22_X1 U793 ( .A1(n97), .A2(\REGISTERS[8][7] ), .B1(n96), .B2(
        \REGISTERS[23][7] ), .ZN(n756) );
  AOI22_X1 U794 ( .A1(n825), .A2(\REGISTERS[16][7] ), .B1(n98), .B2(
        \REGISTERS[1][7] ), .ZN(n755) );
  NAND3_X1 U795 ( .A1(n757), .A2(n756), .A3(n755), .ZN(n758) );
  NOR4_X1 U796 ( .A1(n761), .A2(n760), .A3(n759), .A4(n758), .ZN(n762) );
  NAND4_X1 U797 ( .A1(n765), .A2(n764), .A3(n763), .A4(n762), .ZN(OUT1[7]) );
  AOI22_X1 U798 ( .A1(n71), .A2(\REGISTERS[18][8] ), .B1(n70), .B2(
        \REGISTERS[19][8] ), .ZN(n785) );
  AOI22_X1 U799 ( .A1(n73), .A2(\REGISTERS[20][8] ), .B1(n72), .B2(
        \REGISTERS[21][8] ), .ZN(n784) );
  AOI22_X1 U800 ( .A1(n75), .A2(\REGISTERS[4][8] ), .B1(n74), .B2(
        \REGISTERS[2][8] ), .ZN(n783) );
  AOI22_X1 U801 ( .A1(n77), .A2(\REGISTERS[26][8] ), .B1(n76), .B2(
        \REGISTERS[27][8] ), .ZN(n769) );
  AOI22_X1 U802 ( .A1(n79), .A2(\REGISTERS[28][8] ), .B1(n78), .B2(
        \REGISTERS[29][8] ), .ZN(n768) );
  AOI22_X1 U803 ( .A1(n81), .A2(\REGISTERS[30][8] ), .B1(n80), .B2(
        \REGISTERS[7][8] ), .ZN(n767) );
  AOI22_X1 U804 ( .A1(n83), .A2(\REGISTERS[5][8] ), .B1(n82), .B2(
        \REGISTERS[3][8] ), .ZN(n766) );
  NAND4_X1 U805 ( .A1(n769), .A2(n768), .A3(n767), .A4(n766), .ZN(n781) );
  AOI22_X1 U806 ( .A1(n85), .A2(\REGISTERS[9][8] ), .B1(n84), .B2(
        \REGISTERS[10][8] ), .ZN(n773) );
  AOI22_X1 U807 ( .A1(n87), .A2(\REGISTERS[11][8] ), .B1(n86), .B2(
        \REGISTERS[12][8] ), .ZN(n772) );
  AOI22_X1 U808 ( .A1(n89), .A2(\REGISTERS[13][8] ), .B1(n88), .B2(
        \REGISTERS[14][8] ), .ZN(n771) );
  AOI22_X1 U809 ( .A1(n91), .A2(\REGISTERS[15][8] ), .B1(n90), .B2(
        \REGISTERS[17][8] ), .ZN(n770) );
  NAND4_X1 U810 ( .A1(n773), .A2(n772), .A3(n771), .A4(n770), .ZN(n780) );
  AOI22_X1 U811 ( .A1(n93), .A2(\REGISTERS[31][8] ), .B1(n92), .B2(
        \REGISTERS[22][8] ), .ZN(n774) );
  OAI21_X1 U812 ( .B1(n819), .B2(n68), .A(n774), .ZN(n779) );
  AOI22_X1 U813 ( .A1(n95), .A2(\REGISTERS[24][8] ), .B1(n94), .B2(
        \REGISTERS[25][8] ), .ZN(n777) );
  AOI22_X1 U814 ( .A1(n97), .A2(\REGISTERS[8][8] ), .B1(n96), .B2(
        \REGISTERS[23][8] ), .ZN(n776) );
  AOI22_X1 U815 ( .A1(n825), .A2(\REGISTERS[16][8] ), .B1(n98), .B2(
        \REGISTERS[1][8] ), .ZN(n775) );
  NAND3_X1 U816 ( .A1(n777), .A2(n776), .A3(n775), .ZN(n778) );
  NOR4_X1 U817 ( .A1(n781), .A2(n780), .A3(n779), .A4(n778), .ZN(n782) );
  NAND4_X1 U818 ( .A1(n785), .A2(n784), .A3(n783), .A4(n782), .ZN(OUT1[8]) );
  AOI22_X1 U819 ( .A1(n71), .A2(\REGISTERS[18][9] ), .B1(n70), .B2(
        \REGISTERS[19][9] ), .ZN(n836) );
  AOI22_X1 U820 ( .A1(n73), .A2(\REGISTERS[20][9] ), .B1(n72), .B2(
        \REGISTERS[21][9] ), .ZN(n835) );
  AOI22_X1 U821 ( .A1(n75), .A2(\REGISTERS[4][9] ), .B1(n74), .B2(
        \REGISTERS[2][9] ), .ZN(n834) );
  AOI22_X1 U822 ( .A1(n77), .A2(\REGISTERS[26][9] ), .B1(n76), .B2(
        \REGISTERS[27][9] ), .ZN(n803) );
  AOI22_X1 U823 ( .A1(n79), .A2(\REGISTERS[28][9] ), .B1(n78), .B2(
        \REGISTERS[29][9] ), .ZN(n802) );
  AOI22_X1 U824 ( .A1(n81), .A2(\REGISTERS[30][9] ), .B1(n80), .B2(
        \REGISTERS[7][9] ), .ZN(n801) );
  AOI22_X1 U825 ( .A1(n83), .A2(\REGISTERS[5][9] ), .B1(n82), .B2(
        \REGISTERS[3][9] ), .ZN(n800) );
  NAND4_X1 U826 ( .A1(n803), .A2(n802), .A3(n801), .A4(n800), .ZN(n832) );
  AOI22_X1 U827 ( .A1(n85), .A2(\REGISTERS[9][9] ), .B1(n84), .B2(
        \REGISTERS[10][9] ), .ZN(n815) );
  AOI22_X1 U828 ( .A1(n87), .A2(\REGISTERS[11][9] ), .B1(n86), .B2(
        \REGISTERS[12][9] ), .ZN(n814) );
  AOI22_X1 U829 ( .A1(n89), .A2(\REGISTERS[13][9] ), .B1(n88), .B2(
        \REGISTERS[14][9] ), .ZN(n813) );
  AOI22_X1 U830 ( .A1(n91), .A2(\REGISTERS[15][9] ), .B1(n90), .B2(
        \REGISTERS[17][9] ), .ZN(n812) );
  NAND4_X1 U831 ( .A1(n815), .A2(n814), .A3(n813), .A4(n812), .ZN(n831) );
  AOI22_X1 U832 ( .A1(n93), .A2(\REGISTERS[31][9] ), .B1(n92), .B2(
        \REGISTERS[22][9] ), .ZN(n818) );
  OAI21_X1 U833 ( .B1(n819), .B2(n69), .A(n818), .ZN(n830) );
  AOI22_X1 U834 ( .A1(n95), .A2(\REGISTERS[24][9] ), .B1(n94), .B2(
        \REGISTERS[25][9] ), .ZN(n828) );
  AOI22_X1 U835 ( .A1(n97), .A2(\REGISTERS[8][9] ), .B1(n96), .B2(
        \REGISTERS[23][9] ), .ZN(n827) );
  AOI22_X1 U836 ( .A1(n825), .A2(\REGISTERS[16][9] ), .B1(n98), .B2(
        \REGISTERS[1][9] ), .ZN(n826) );
  NAND3_X1 U837 ( .A1(n828), .A2(n827), .A3(n826), .ZN(n829) );
  NOR4_X1 U838 ( .A1(n832), .A2(n831), .A3(n830), .A4(n829), .ZN(n833) );
  NAND4_X1 U839 ( .A1(n836), .A2(n835), .A3(n834), .A4(n833), .ZN(OUT1[9]) );
  INV_X1 U840 ( .A(ADD_RD2[2]), .ZN(n840) );
  NAND2_X1 U841 ( .A1(ADD_RD2[1]), .A2(n840), .ZN(n850) );
  INV_X1 U842 ( .A(ADD_RD2[0]), .ZN(n869) );
  INV_X1 U843 ( .A(ADD_RD2[3]), .ZN(n837) );
  NAND3_X1 U844 ( .A1(ADD_RD2[4]), .A2(n869), .A3(n837), .ZN(n860) );
  NOR2_X1 U845 ( .A1(n850), .A2(n860), .ZN(n1482) );
  NAND3_X1 U846 ( .A1(ADD_RD2[4]), .A2(ADD_RD2[0]), .A3(n837), .ZN(n865) );
  NOR2_X1 U847 ( .A1(n850), .A2(n865), .ZN(n1481) );
  AOI22_X1 U848 ( .A1(\REGISTERS[18][0] ), .A2(n100), .B1(\REGISTERS[19][0] ), 
        .B2(n99), .ZN(n880) );
  INV_X1 U849 ( .A(ADD_RD2[1]), .ZN(n841) );
  NAND2_X1 U850 ( .A1(ADD_RD2[2]), .A2(n841), .ZN(n851) );
  NOR2_X1 U851 ( .A1(n851), .A2(n860), .ZN(n1484) );
  NOR2_X1 U852 ( .A1(n851), .A2(n865), .ZN(n1483) );
  AOI22_X1 U853 ( .A1(\REGISTERS[20][0] ), .A2(n102), .B1(\REGISTERS[21][0] ), 
        .B2(n101), .ZN(n879) );
  NOR3_X1 U854 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[4]), .A3(ADD_RD2[3]), .ZN(n858)
         );
  NAND2_X1 U855 ( .A1(n841), .A2(n840), .ZN(n868) );
  NOR3_X1 U856 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[3]), .A3(n868), .ZN(n867) );
  INV_X1 U857 ( .A(ADD_RD2[4]), .ZN(n848) );
  NAND2_X1 U858 ( .A1(n867), .A2(n848), .ZN(n838) );
  NAND2_X1 U859 ( .A1(n858), .A2(n838), .ZN(n839) );
  NOR2_X1 U860 ( .A1(ADD_RD2[1]), .A2(n839), .ZN(n1486) );
  NOR2_X1 U861 ( .A1(ADD_RD2[2]), .A2(n839), .ZN(n1485) );
  AOI22_X1 U862 ( .A1(\REGISTERS[4][0] ), .A2(n104), .B1(\REGISTERS[2][0] ), 
        .B2(n103), .ZN(n878) );
  NAND3_X1 U863 ( .A1(ADD_RD2[4]), .A2(ADD_RD2[3]), .A3(n869), .ZN(n862) );
  NOR2_X1 U864 ( .A1(n862), .A2(n850), .ZN(n1488) );
  NAND3_X1 U865 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[4]), .A3(ADD_RD2[3]), .ZN(n863)
         );
  NOR2_X1 U866 ( .A1(n850), .A2(n863), .ZN(n1487) );
  AOI22_X1 U867 ( .A1(\REGISTERS[26][0] ), .A2(n106), .B1(\REGISTERS[27][0] ), 
        .B2(n105), .ZN(n847) );
  NOR2_X1 U868 ( .A1(n862), .A2(n851), .ZN(n1490) );
  NOR2_X1 U869 ( .A1(n863), .A2(n851), .ZN(n1489) );
  AOI22_X1 U870 ( .A1(\REGISTERS[28][0] ), .A2(n108), .B1(\REGISTERS[29][0] ), 
        .B2(n107), .ZN(n846) );
  NOR2_X1 U871 ( .A1(n841), .A2(n840), .ZN(n859) );
  INV_X1 U872 ( .A(n859), .ZN(n866) );
  NOR2_X1 U873 ( .A1(n862), .A2(n866), .ZN(n1492) );
  NOR2_X1 U874 ( .A1(ADD_RD2[4]), .A2(ADD_RD2[3]), .ZN(n842) );
  NAND2_X1 U875 ( .A1(ADD_RD2[0]), .A2(n842), .ZN(n843) );
  NOR2_X1 U876 ( .A1(n866), .A2(n843), .ZN(n1491) );
  AOI22_X1 U877 ( .A1(\REGISTERS[30][0] ), .A2(n110), .B1(\REGISTERS[7][0] ), 
        .B2(n109), .ZN(n845) );
  NOR2_X1 U878 ( .A1(n851), .A2(n843), .ZN(n1494) );
  NOR2_X1 U879 ( .A1(n850), .A2(n843), .ZN(n1493) );
  AOI22_X1 U880 ( .A1(\REGISTERS[5][0] ), .A2(n112), .B1(\REGISTERS[3][0] ), 
        .B2(n111), .ZN(n844) );
  NAND4_X1 U881 ( .A1(n847), .A2(n846), .A3(n845), .A4(n844), .ZN(n876) );
  NAND2_X1 U882 ( .A1(n848), .A2(ADD_RD2[3]), .ZN(n864) );
  INV_X1 U883 ( .A(n864), .ZN(n849) );
  NAND2_X1 U884 ( .A1(ADD_RD2[0]), .A2(n849), .ZN(n853) );
  NOR2_X1 U885 ( .A1(n868), .A2(n853), .ZN(n1500) );
  NAND2_X1 U886 ( .A1(n849), .A2(n869), .ZN(n852) );
  NOR2_X1 U887 ( .A1(n850), .A2(n852), .ZN(n1499) );
  AOI22_X1 U888 ( .A1(\REGISTERS[9][0] ), .A2(n114), .B1(\REGISTERS[10][0] ), 
        .B2(n113), .ZN(n857) );
  NOR2_X1 U889 ( .A1(n850), .A2(n853), .ZN(n1502) );
  NOR2_X1 U890 ( .A1(n851), .A2(n852), .ZN(n1501) );
  AOI22_X1 U891 ( .A1(\REGISTERS[11][0] ), .A2(n116), .B1(\REGISTERS[12][0] ), 
        .B2(n115), .ZN(n856) );
  NOR2_X1 U892 ( .A1(n851), .A2(n853), .ZN(n1504) );
  NOR2_X1 U893 ( .A1(n866), .A2(n852), .ZN(n1503) );
  AOI22_X1 U894 ( .A1(\REGISTERS[13][0] ), .A2(n118), .B1(\REGISTERS[14][0] ), 
        .B2(n117), .ZN(n855) );
  NOR2_X1 U895 ( .A1(n866), .A2(n853), .ZN(n1506) );
  NOR2_X1 U896 ( .A1(n868), .A2(n865), .ZN(n1505) );
  AOI22_X1 U897 ( .A1(\REGISTERS[15][0] ), .A2(n120), .B1(\REGISTERS[17][0] ), 
        .B2(n119), .ZN(n854) );
  NAND4_X1 U898 ( .A1(n857), .A2(n856), .A3(n855), .A4(n854), .ZN(n875) );
  NOR2_X1 U899 ( .A1(n863), .A2(n866), .ZN(n1512) );
  NOR2_X1 U900 ( .A1(n866), .A2(n860), .ZN(n1511) );
  AOI22_X1 U901 ( .A1(\REGISTERS[31][0] ), .A2(n122), .B1(\REGISTERS[22][0] ), 
        .B2(n121), .ZN(n861) );
  OAI21_X1 U902 ( .B1(n38), .B2(n1514), .A(n861), .ZN(n874) );
  NOR2_X1 U903 ( .A1(n862), .A2(n868), .ZN(n1516) );
  NOR2_X1 U904 ( .A1(n863), .A2(n868), .ZN(n1515) );
  AOI22_X1 U905 ( .A1(\REGISTERS[24][0] ), .A2(n124), .B1(\REGISTERS[25][0] ), 
        .B2(n123), .ZN(n872) );
  NOR3_X1 U906 ( .A1(ADD_RD2[0]), .A2(n868), .A3(n864), .ZN(n1518) );
  NOR2_X1 U907 ( .A1(n866), .A2(n865), .ZN(n1517) );
  AOI22_X1 U908 ( .A1(\REGISTERS[8][0] ), .A2(n36), .B1(\REGISTERS[23][0] ), 
        .B2(n125), .ZN(n871) );
  NOR4_X1 U909 ( .A1(ADD_RD2[3]), .A2(ADD_RD2[4]), .A3(n869), .A4(n868), .ZN(
        n1519) );
  AOI22_X1 U910 ( .A1(\REGISTERS[16][0] ), .A2(n1520), .B1(\REGISTERS[1][0] ), 
        .B2(n37), .ZN(n870) );
  NAND3_X1 U911 ( .A1(n872), .A2(n871), .A3(n870), .ZN(n873) );
  NOR4_X1 U912 ( .A1(n876), .A2(n875), .A3(n874), .A4(n873), .ZN(n877) );
  NAND4_X1 U913 ( .A1(n880), .A2(n879), .A3(n878), .A4(n877), .ZN(OUT2[0]) );
  AOI22_X1 U914 ( .A1(\REGISTERS[18][10] ), .A2(n100), .B1(\REGISTERS[19][10] ), .B2(n99), .ZN(n900) );
  AOI22_X1 U915 ( .A1(\REGISTERS[20][10] ), .A2(n102), .B1(\REGISTERS[21][10] ), .B2(n101), .ZN(n899) );
  AOI22_X1 U916 ( .A1(\REGISTERS[4][10] ), .A2(n104), .B1(\REGISTERS[2][10] ), 
        .B2(n103), .ZN(n898) );
  AOI22_X1 U917 ( .A1(\REGISTERS[26][10] ), .A2(n106), .B1(\REGISTERS[27][10] ), .B2(n105), .ZN(n884) );
  AOI22_X1 U918 ( .A1(\REGISTERS[28][10] ), .A2(n108), .B1(\REGISTERS[29][10] ), .B2(n107), .ZN(n883) );
  AOI22_X1 U919 ( .A1(\REGISTERS[30][10] ), .A2(n110), .B1(\REGISTERS[7][10] ), 
        .B2(n109), .ZN(n882) );
  AOI22_X1 U920 ( .A1(\REGISTERS[5][10] ), .A2(n112), .B1(\REGISTERS[3][10] ), 
        .B2(n111), .ZN(n881) );
  NAND4_X1 U921 ( .A1(n884), .A2(n883), .A3(n882), .A4(n881), .ZN(n896) );
  AOI22_X1 U922 ( .A1(\REGISTERS[9][10] ), .A2(n114), .B1(\REGISTERS[10][10] ), 
        .B2(n113), .ZN(n888) );
  AOI22_X1 U923 ( .A1(\REGISTERS[11][10] ), .A2(n116), .B1(\REGISTERS[12][10] ), .B2(n115), .ZN(n887) );
  AOI22_X1 U924 ( .A1(\REGISTERS[13][10] ), .A2(n118), .B1(\REGISTERS[14][10] ), .B2(n117), .ZN(n886) );
  AOI22_X1 U925 ( .A1(\REGISTERS[15][10] ), .A2(n120), .B1(\REGISTERS[17][10] ), .B2(n119), .ZN(n885) );
  NAND4_X1 U926 ( .A1(n888), .A2(n887), .A3(n886), .A4(n885), .ZN(n895) );
  AOI22_X1 U927 ( .A1(\REGISTERS[31][10] ), .A2(n122), .B1(\REGISTERS[22][10] ), .B2(n121), .ZN(n889) );
  OAI21_X1 U928 ( .B1(n39), .B2(n1514), .A(n889), .ZN(n894) );
  AOI22_X1 U929 ( .A1(\REGISTERS[24][10] ), .A2(n124), .B1(\REGISTERS[25][10] ), .B2(n123), .ZN(n892) );
  AOI22_X1 U930 ( .A1(\REGISTERS[8][10] ), .A2(n36), .B1(\REGISTERS[23][10] ), 
        .B2(n125), .ZN(n891) );
  AOI22_X1 U931 ( .A1(\REGISTERS[16][10] ), .A2(n1520), .B1(\REGISTERS[1][10] ), .B2(n37), .ZN(n890) );
  NAND3_X1 U932 ( .A1(n892), .A2(n891), .A3(n890), .ZN(n893) );
  NOR4_X1 U933 ( .A1(n896), .A2(n895), .A3(n894), .A4(n893), .ZN(n897) );
  NAND4_X1 U934 ( .A1(n900), .A2(n899), .A3(n898), .A4(n897), .ZN(OUT2[10]) );
  AOI22_X1 U935 ( .A1(\REGISTERS[18][11] ), .A2(n100), .B1(\REGISTERS[19][11] ), .B2(n99), .ZN(n920) );
  AOI22_X1 U936 ( .A1(\REGISTERS[20][11] ), .A2(n102), .B1(\REGISTERS[21][11] ), .B2(n101), .ZN(n919) );
  AOI22_X1 U937 ( .A1(\REGISTERS[4][11] ), .A2(n104), .B1(\REGISTERS[2][11] ), 
        .B2(n103), .ZN(n918) );
  AOI22_X1 U938 ( .A1(\REGISTERS[26][11] ), .A2(n106), .B1(\REGISTERS[27][11] ), .B2(n105), .ZN(n904) );
  AOI22_X1 U939 ( .A1(\REGISTERS[28][11] ), .A2(n108), .B1(\REGISTERS[29][11] ), .B2(n107), .ZN(n903) );
  AOI22_X1 U940 ( .A1(\REGISTERS[30][11] ), .A2(n110), .B1(\REGISTERS[7][11] ), 
        .B2(n109), .ZN(n902) );
  AOI22_X1 U941 ( .A1(\REGISTERS[5][11] ), .A2(n112), .B1(\REGISTERS[3][11] ), 
        .B2(n111), .ZN(n901) );
  NAND4_X1 U942 ( .A1(n904), .A2(n903), .A3(n902), .A4(n901), .ZN(n916) );
  AOI22_X1 U943 ( .A1(\REGISTERS[9][11] ), .A2(n114), .B1(\REGISTERS[10][11] ), 
        .B2(n113), .ZN(n908) );
  AOI22_X1 U944 ( .A1(\REGISTERS[11][11] ), .A2(n116), .B1(\REGISTERS[12][11] ), .B2(n115), .ZN(n907) );
  AOI22_X1 U945 ( .A1(\REGISTERS[13][11] ), .A2(n118), .B1(\REGISTERS[14][11] ), .B2(n117), .ZN(n906) );
  AOI22_X1 U946 ( .A1(\REGISTERS[15][11] ), .A2(n120), .B1(\REGISTERS[17][11] ), .B2(n119), .ZN(n905) );
  NAND4_X1 U947 ( .A1(n908), .A2(n907), .A3(n906), .A4(n905), .ZN(n915) );
  AOI22_X1 U948 ( .A1(\REGISTERS[31][11] ), .A2(n122), .B1(\REGISTERS[22][11] ), .B2(n121), .ZN(n909) );
  OAI21_X1 U949 ( .B1(n40), .B2(n1514), .A(n909), .ZN(n914) );
  AOI22_X1 U950 ( .A1(\REGISTERS[24][11] ), .A2(n124), .B1(\REGISTERS[25][11] ), .B2(n123), .ZN(n912) );
  AOI22_X1 U951 ( .A1(\REGISTERS[8][11] ), .A2(n36), .B1(\REGISTERS[23][11] ), 
        .B2(n125), .ZN(n911) );
  AOI22_X1 U952 ( .A1(\REGISTERS[16][11] ), .A2(n1520), .B1(\REGISTERS[1][11] ), .B2(n37), .ZN(n910) );
  NAND3_X1 U953 ( .A1(n912), .A2(n911), .A3(n910), .ZN(n913) );
  NOR4_X1 U954 ( .A1(n916), .A2(n915), .A3(n914), .A4(n913), .ZN(n917) );
  NAND4_X1 U955 ( .A1(n920), .A2(n919), .A3(n918), .A4(n917), .ZN(OUT2[11]) );
  AOI22_X1 U956 ( .A1(\REGISTERS[18][12] ), .A2(n100), .B1(\REGISTERS[19][12] ), .B2(n99), .ZN(n940) );
  AOI22_X1 U957 ( .A1(\REGISTERS[20][12] ), .A2(n102), .B1(\REGISTERS[21][12] ), .B2(n101), .ZN(n939) );
  AOI22_X1 U958 ( .A1(\REGISTERS[4][12] ), .A2(n104), .B1(\REGISTERS[2][12] ), 
        .B2(n103), .ZN(n938) );
  AOI22_X1 U959 ( .A1(\REGISTERS[26][12] ), .A2(n106), .B1(\REGISTERS[27][12] ), .B2(n105), .ZN(n924) );
  AOI22_X1 U960 ( .A1(\REGISTERS[28][12] ), .A2(n108), .B1(\REGISTERS[29][12] ), .B2(n107), .ZN(n923) );
  AOI22_X1 U961 ( .A1(\REGISTERS[30][12] ), .A2(n110), .B1(\REGISTERS[7][12] ), 
        .B2(n109), .ZN(n922) );
  AOI22_X1 U962 ( .A1(\REGISTERS[5][12] ), .A2(n112), .B1(\REGISTERS[3][12] ), 
        .B2(n111), .ZN(n921) );
  NAND4_X1 U963 ( .A1(n924), .A2(n923), .A3(n922), .A4(n921), .ZN(n936) );
  AOI22_X1 U964 ( .A1(\REGISTERS[9][12] ), .A2(n114), .B1(\REGISTERS[10][12] ), 
        .B2(n113), .ZN(n928) );
  AOI22_X1 U965 ( .A1(\REGISTERS[11][12] ), .A2(n116), .B1(\REGISTERS[12][12] ), .B2(n115), .ZN(n927) );
  AOI22_X1 U966 ( .A1(\REGISTERS[13][12] ), .A2(n118), .B1(\REGISTERS[14][12] ), .B2(n117), .ZN(n926) );
  AOI22_X1 U967 ( .A1(\REGISTERS[15][12] ), .A2(n120), .B1(\REGISTERS[17][12] ), .B2(n119), .ZN(n925) );
  NAND4_X1 U968 ( .A1(n928), .A2(n927), .A3(n926), .A4(n925), .ZN(n935) );
  AOI22_X1 U969 ( .A1(\REGISTERS[31][12] ), .A2(n122), .B1(\REGISTERS[22][12] ), .B2(n121), .ZN(n929) );
  OAI21_X1 U970 ( .B1(n41), .B2(n1514), .A(n929), .ZN(n934) );
  AOI22_X1 U971 ( .A1(\REGISTERS[24][12] ), .A2(n124), .B1(\REGISTERS[25][12] ), .B2(n123), .ZN(n932) );
  AOI22_X1 U972 ( .A1(\REGISTERS[8][12] ), .A2(n36), .B1(\REGISTERS[23][12] ), 
        .B2(n125), .ZN(n931) );
  AOI22_X1 U973 ( .A1(\REGISTERS[16][12] ), .A2(n1520), .B1(\REGISTERS[1][12] ), .B2(n37), .ZN(n930) );
  NAND3_X1 U974 ( .A1(n932), .A2(n931), .A3(n930), .ZN(n933) );
  NOR4_X1 U975 ( .A1(n936), .A2(n935), .A3(n934), .A4(n933), .ZN(n937) );
  NAND4_X1 U976 ( .A1(n940), .A2(n939), .A3(n938), .A4(n937), .ZN(OUT2[12]) );
  AOI22_X1 U977 ( .A1(\REGISTERS[18][13] ), .A2(n100), .B1(\REGISTERS[19][13] ), .B2(n99), .ZN(n960) );
  AOI22_X1 U978 ( .A1(\REGISTERS[20][13] ), .A2(n102), .B1(\REGISTERS[21][13] ), .B2(n101), .ZN(n959) );
  AOI22_X1 U979 ( .A1(\REGISTERS[4][13] ), .A2(n104), .B1(\REGISTERS[2][13] ), 
        .B2(n103), .ZN(n958) );
  AOI22_X1 U980 ( .A1(\REGISTERS[26][13] ), .A2(n106), .B1(\REGISTERS[27][13] ), .B2(n105), .ZN(n944) );
  AOI22_X1 U981 ( .A1(\REGISTERS[28][13] ), .A2(n108), .B1(\REGISTERS[29][13] ), .B2(n107), .ZN(n943) );
  AOI22_X1 U982 ( .A1(\REGISTERS[30][13] ), .A2(n110), .B1(\REGISTERS[7][13] ), 
        .B2(n109), .ZN(n942) );
  AOI22_X1 U983 ( .A1(\REGISTERS[5][13] ), .A2(n112), .B1(\REGISTERS[3][13] ), 
        .B2(n111), .ZN(n941) );
  NAND4_X1 U984 ( .A1(n944), .A2(n943), .A3(n942), .A4(n941), .ZN(n956) );
  AOI22_X1 U985 ( .A1(\REGISTERS[9][13] ), .A2(n114), .B1(\REGISTERS[10][13] ), 
        .B2(n113), .ZN(n948) );
  AOI22_X1 U986 ( .A1(\REGISTERS[11][13] ), .A2(n116), .B1(\REGISTERS[12][13] ), .B2(n115), .ZN(n947) );
  AOI22_X1 U987 ( .A1(\REGISTERS[13][13] ), .A2(n118), .B1(\REGISTERS[14][13] ), .B2(n117), .ZN(n946) );
  AOI22_X1 U988 ( .A1(\REGISTERS[15][13] ), .A2(n120), .B1(\REGISTERS[17][13] ), .B2(n119), .ZN(n945) );
  NAND4_X1 U989 ( .A1(n948), .A2(n947), .A3(n946), .A4(n945), .ZN(n955) );
  AOI22_X1 U990 ( .A1(\REGISTERS[31][13] ), .A2(n122), .B1(\REGISTERS[22][13] ), .B2(n121), .ZN(n949) );
  OAI21_X1 U991 ( .B1(n42), .B2(n1514), .A(n949), .ZN(n954) );
  AOI22_X1 U992 ( .A1(\REGISTERS[24][13] ), .A2(n124), .B1(\REGISTERS[25][13] ), .B2(n123), .ZN(n952) );
  AOI22_X1 U993 ( .A1(\REGISTERS[8][13] ), .A2(n36), .B1(\REGISTERS[23][13] ), 
        .B2(n125), .ZN(n951) );
  AOI22_X1 U994 ( .A1(\REGISTERS[16][13] ), .A2(n1520), .B1(\REGISTERS[1][13] ), .B2(n37), .ZN(n950) );
  NAND3_X1 U995 ( .A1(n952), .A2(n951), .A3(n950), .ZN(n953) );
  NOR4_X1 U996 ( .A1(n956), .A2(n955), .A3(n954), .A4(n953), .ZN(n957) );
  NAND4_X1 U997 ( .A1(n960), .A2(n959), .A3(n958), .A4(n957), .ZN(OUT2[13]) );
  AOI22_X1 U998 ( .A1(\REGISTERS[18][14] ), .A2(n100), .B1(\REGISTERS[19][14] ), .B2(n99), .ZN(n980) );
  AOI22_X1 U999 ( .A1(\REGISTERS[20][14] ), .A2(n102), .B1(\REGISTERS[21][14] ), .B2(n101), .ZN(n979) );
  AOI22_X1 U1000 ( .A1(\REGISTERS[4][14] ), .A2(n104), .B1(\REGISTERS[2][14] ), 
        .B2(n103), .ZN(n978) );
  AOI22_X1 U1001 ( .A1(\REGISTERS[26][14] ), .A2(n106), .B1(
        \REGISTERS[27][14] ), .B2(n105), .ZN(n964) );
  AOI22_X1 U1002 ( .A1(\REGISTERS[28][14] ), .A2(n108), .B1(
        \REGISTERS[29][14] ), .B2(n107), .ZN(n963) );
  AOI22_X1 U1003 ( .A1(\REGISTERS[30][14] ), .A2(n110), .B1(\REGISTERS[7][14] ), .B2(n109), .ZN(n962) );
  AOI22_X1 U1004 ( .A1(\REGISTERS[5][14] ), .A2(n112), .B1(\REGISTERS[3][14] ), 
        .B2(n111), .ZN(n961) );
  NAND4_X1 U1005 ( .A1(n964), .A2(n963), .A3(n962), .A4(n961), .ZN(n976) );
  AOI22_X1 U1006 ( .A1(\REGISTERS[9][14] ), .A2(n114), .B1(\REGISTERS[10][14] ), .B2(n113), .ZN(n968) );
  AOI22_X1 U1007 ( .A1(\REGISTERS[11][14] ), .A2(n116), .B1(
        \REGISTERS[12][14] ), .B2(n115), .ZN(n967) );
  AOI22_X1 U1008 ( .A1(\REGISTERS[13][14] ), .A2(n118), .B1(
        \REGISTERS[14][14] ), .B2(n117), .ZN(n966) );
  AOI22_X1 U1009 ( .A1(\REGISTERS[15][14] ), .A2(n120), .B1(
        \REGISTERS[17][14] ), .B2(n119), .ZN(n965) );
  NAND4_X1 U1010 ( .A1(n968), .A2(n967), .A3(n966), .A4(n965), .ZN(n975) );
  AOI22_X1 U1011 ( .A1(\REGISTERS[31][14] ), .A2(n122), .B1(
        \REGISTERS[22][14] ), .B2(n121), .ZN(n969) );
  OAI21_X1 U1012 ( .B1(n43), .B2(n1514), .A(n969), .ZN(n974) );
  AOI22_X1 U1013 ( .A1(\REGISTERS[24][14] ), .A2(n124), .B1(
        \REGISTERS[25][14] ), .B2(n123), .ZN(n972) );
  AOI22_X1 U1014 ( .A1(\REGISTERS[8][14] ), .A2(n36), .B1(\REGISTERS[23][14] ), 
        .B2(n125), .ZN(n971) );
  AOI22_X1 U1015 ( .A1(\REGISTERS[16][14] ), .A2(n1520), .B1(
        \REGISTERS[1][14] ), .B2(n37), .ZN(n970) );
  NAND3_X1 U1016 ( .A1(n972), .A2(n971), .A3(n970), .ZN(n973) );
  NOR4_X1 U1017 ( .A1(n976), .A2(n975), .A3(n974), .A4(n973), .ZN(n977) );
  NAND4_X1 U1018 ( .A1(n980), .A2(n979), .A3(n978), .A4(n977), .ZN(OUT2[14])
         );
  AOI22_X1 U1019 ( .A1(\REGISTERS[18][15] ), .A2(n100), .B1(
        \REGISTERS[19][15] ), .B2(n99), .ZN(n1000) );
  AOI22_X1 U1020 ( .A1(\REGISTERS[20][15] ), .A2(n102), .B1(
        \REGISTERS[21][15] ), .B2(n101), .ZN(n999) );
  AOI22_X1 U1021 ( .A1(\REGISTERS[4][15] ), .A2(n104), .B1(\REGISTERS[2][15] ), 
        .B2(n103), .ZN(n998) );
  AOI22_X1 U1022 ( .A1(\REGISTERS[26][15] ), .A2(n106), .B1(
        \REGISTERS[27][15] ), .B2(n105), .ZN(n984) );
  AOI22_X1 U1023 ( .A1(\REGISTERS[28][15] ), .A2(n108), .B1(
        \REGISTERS[29][15] ), .B2(n107), .ZN(n983) );
  AOI22_X1 U1024 ( .A1(\REGISTERS[30][15] ), .A2(n110), .B1(\REGISTERS[7][15] ), .B2(n109), .ZN(n982) );
  AOI22_X1 U1025 ( .A1(\REGISTERS[5][15] ), .A2(n112), .B1(\REGISTERS[3][15] ), 
        .B2(n111), .ZN(n981) );
  NAND4_X1 U1026 ( .A1(n984), .A2(n983), .A3(n982), .A4(n981), .ZN(n996) );
  AOI22_X1 U1027 ( .A1(\REGISTERS[9][15] ), .A2(n114), .B1(\REGISTERS[10][15] ), .B2(n113), .ZN(n988) );
  AOI22_X1 U1028 ( .A1(\REGISTERS[11][15] ), .A2(n116), .B1(
        \REGISTERS[12][15] ), .B2(n115), .ZN(n987) );
  AOI22_X1 U1029 ( .A1(\REGISTERS[13][15] ), .A2(n118), .B1(
        \REGISTERS[14][15] ), .B2(n117), .ZN(n986) );
  AOI22_X1 U1030 ( .A1(\REGISTERS[15][15] ), .A2(n120), .B1(
        \REGISTERS[17][15] ), .B2(n119), .ZN(n985) );
  NAND4_X1 U1031 ( .A1(n988), .A2(n987), .A3(n986), .A4(n985), .ZN(n995) );
  AOI22_X1 U1032 ( .A1(\REGISTERS[31][15] ), .A2(n122), .B1(
        \REGISTERS[22][15] ), .B2(n121), .ZN(n989) );
  OAI21_X1 U1033 ( .B1(n44), .B2(n1514), .A(n989), .ZN(n994) );
  AOI22_X1 U1034 ( .A1(\REGISTERS[24][15] ), .A2(n124), .B1(
        \REGISTERS[25][15] ), .B2(n123), .ZN(n992) );
  AOI22_X1 U1035 ( .A1(\REGISTERS[8][15] ), .A2(n36), .B1(\REGISTERS[23][15] ), 
        .B2(n125), .ZN(n991) );
  AOI22_X1 U1036 ( .A1(\REGISTERS[16][15] ), .A2(n1520), .B1(
        \REGISTERS[1][15] ), .B2(n37), .ZN(n990) );
  NAND3_X1 U1037 ( .A1(n992), .A2(n991), .A3(n990), .ZN(n993) );
  NOR4_X1 U1038 ( .A1(n996), .A2(n995), .A3(n994), .A4(n993), .ZN(n997) );
  NAND4_X1 U1039 ( .A1(n1000), .A2(n999), .A3(n998), .A4(n997), .ZN(OUT2[15])
         );
  AOI22_X1 U1040 ( .A1(\REGISTERS[18][16] ), .A2(n1482), .B1(
        \REGISTERS[19][16] ), .B2(n99), .ZN(n1020) );
  AOI22_X1 U1041 ( .A1(\REGISTERS[20][16] ), .A2(n1484), .B1(
        \REGISTERS[21][16] ), .B2(n101), .ZN(n1019) );
  AOI22_X1 U1042 ( .A1(\REGISTERS[4][16] ), .A2(n1486), .B1(\REGISTERS[2][16] ), .B2(n103), .ZN(n1018) );
  AOI22_X1 U1043 ( .A1(\REGISTERS[26][16] ), .A2(n106), .B1(
        \REGISTERS[27][16] ), .B2(n105), .ZN(n1004) );
  AOI22_X1 U1044 ( .A1(\REGISTERS[28][16] ), .A2(n108), .B1(
        \REGISTERS[29][16] ), .B2(n107), .ZN(n1003) );
  AOI22_X1 U1045 ( .A1(\REGISTERS[30][16] ), .A2(n110), .B1(\REGISTERS[7][16] ), .B2(n109), .ZN(n1002) );
  AOI22_X1 U1046 ( .A1(\REGISTERS[5][16] ), .A2(n112), .B1(\REGISTERS[3][16] ), 
        .B2(n111), .ZN(n1001) );
  NAND4_X1 U1047 ( .A1(n1004), .A2(n1003), .A3(n1002), .A4(n1001), .ZN(n1016)
         );
  AOI22_X1 U1048 ( .A1(\REGISTERS[9][16] ), .A2(n114), .B1(\REGISTERS[10][16] ), .B2(n113), .ZN(n1008) );
  AOI22_X1 U1049 ( .A1(\REGISTERS[11][16] ), .A2(n116), .B1(
        \REGISTERS[12][16] ), .B2(n115), .ZN(n1007) );
  AOI22_X1 U1050 ( .A1(\REGISTERS[13][16] ), .A2(n118), .B1(
        \REGISTERS[14][16] ), .B2(n117), .ZN(n1006) );
  AOI22_X1 U1051 ( .A1(\REGISTERS[15][16] ), .A2(n120), .B1(
        \REGISTERS[17][16] ), .B2(n119), .ZN(n1005) );
  NAND4_X1 U1052 ( .A1(n1008), .A2(n1007), .A3(n1006), .A4(n1005), .ZN(n1015)
         );
  AOI22_X1 U1053 ( .A1(\REGISTERS[31][16] ), .A2(n122), .B1(
        \REGISTERS[22][16] ), .B2(n121), .ZN(n1009) );
  OAI21_X1 U1054 ( .B1(n45), .B2(n1514), .A(n1009), .ZN(n1014) );
  AOI22_X1 U1055 ( .A1(\REGISTERS[24][16] ), .A2(n124), .B1(
        \REGISTERS[25][16] ), .B2(n123), .ZN(n1012) );
  AOI22_X1 U1056 ( .A1(\REGISTERS[8][16] ), .A2(n36), .B1(\REGISTERS[23][16] ), 
        .B2(n125), .ZN(n1011) );
  AOI22_X1 U1057 ( .A1(\REGISTERS[16][16] ), .A2(n1520), .B1(
        \REGISTERS[1][16] ), .B2(n37), .ZN(n1010) );
  NAND3_X1 U1058 ( .A1(n1012), .A2(n1011), .A3(n1010), .ZN(n1013) );
  NOR4_X1 U1059 ( .A1(n1016), .A2(n1015), .A3(n1014), .A4(n1013), .ZN(n1017)
         );
  NAND4_X1 U1060 ( .A1(n1020), .A2(n1019), .A3(n1018), .A4(n1017), .ZN(
        OUT2[16]) );
  AOI22_X1 U1061 ( .A1(\REGISTERS[18][17] ), .A2(n1482), .B1(
        \REGISTERS[19][17] ), .B2(n99), .ZN(n1040) );
  AOI22_X1 U1062 ( .A1(\REGISTERS[20][17] ), .A2(n1484), .B1(
        \REGISTERS[21][17] ), .B2(n101), .ZN(n1039) );
  AOI22_X1 U1063 ( .A1(\REGISTERS[4][17] ), .A2(n1486), .B1(\REGISTERS[2][17] ), .B2(n103), .ZN(n1038) );
  AOI22_X1 U1064 ( .A1(\REGISTERS[26][17] ), .A2(n106), .B1(
        \REGISTERS[27][17] ), .B2(n1487), .ZN(n1024) );
  AOI22_X1 U1065 ( .A1(\REGISTERS[28][17] ), .A2(n108), .B1(
        \REGISTERS[29][17] ), .B2(n1489), .ZN(n1023) );
  AOI22_X1 U1066 ( .A1(\REGISTERS[30][17] ), .A2(n110), .B1(\REGISTERS[7][17] ), .B2(n1491), .ZN(n1022) );
  AOI22_X1 U1067 ( .A1(\REGISTERS[5][17] ), .A2(n112), .B1(\REGISTERS[3][17] ), 
        .B2(n1493), .ZN(n1021) );
  NAND4_X1 U1068 ( .A1(n1024), .A2(n1023), .A3(n1022), .A4(n1021), .ZN(n1036)
         );
  AOI22_X1 U1069 ( .A1(\REGISTERS[9][17] ), .A2(n114), .B1(\REGISTERS[10][17] ), .B2(n113), .ZN(n1028) );
  AOI22_X1 U1070 ( .A1(\REGISTERS[11][17] ), .A2(n116), .B1(
        \REGISTERS[12][17] ), .B2(n115), .ZN(n1027) );
  AOI22_X1 U1071 ( .A1(\REGISTERS[13][17] ), .A2(n118), .B1(
        \REGISTERS[14][17] ), .B2(n117), .ZN(n1026) );
  AOI22_X1 U1072 ( .A1(\REGISTERS[15][17] ), .A2(n120), .B1(
        \REGISTERS[17][17] ), .B2(n119), .ZN(n1025) );
  NAND4_X1 U1073 ( .A1(n1028), .A2(n1027), .A3(n1026), .A4(n1025), .ZN(n1035)
         );
  AOI22_X1 U1074 ( .A1(\REGISTERS[31][17] ), .A2(n122), .B1(
        \REGISTERS[22][17] ), .B2(n121), .ZN(n1029) );
  OAI21_X1 U1075 ( .B1(n46), .B2(n1514), .A(n1029), .ZN(n1034) );
  AOI22_X1 U1076 ( .A1(\REGISTERS[24][17] ), .A2(n124), .B1(
        \REGISTERS[25][17] ), .B2(n1515), .ZN(n1032) );
  AOI22_X1 U1077 ( .A1(\REGISTERS[8][17] ), .A2(n36), .B1(\REGISTERS[23][17] ), 
        .B2(n125), .ZN(n1031) );
  AOI22_X1 U1078 ( .A1(\REGISTERS[16][17] ), .A2(n1520), .B1(
        \REGISTERS[1][17] ), .B2(n37), .ZN(n1030) );
  NAND3_X1 U1079 ( .A1(n1032), .A2(n1031), .A3(n1030), .ZN(n1033) );
  NOR4_X1 U1080 ( .A1(n1036), .A2(n1035), .A3(n1034), .A4(n1033), .ZN(n1037)
         );
  NAND4_X1 U1081 ( .A1(n1040), .A2(n1039), .A3(n1038), .A4(n1037), .ZN(
        OUT2[17]) );
  AOI22_X1 U1082 ( .A1(\REGISTERS[18][18] ), .A2(n100), .B1(
        \REGISTERS[19][18] ), .B2(n1481), .ZN(n1060) );
  AOI22_X1 U1083 ( .A1(\REGISTERS[20][18] ), .A2(n102), .B1(
        \REGISTERS[21][18] ), .B2(n1483), .ZN(n1059) );
  AOI22_X1 U1084 ( .A1(\REGISTERS[4][18] ), .A2(n104), .B1(\REGISTERS[2][18] ), 
        .B2(n1485), .ZN(n1058) );
  AOI22_X1 U1085 ( .A1(\REGISTERS[26][18] ), .A2(n106), .B1(
        \REGISTERS[27][18] ), .B2(n1487), .ZN(n1044) );
  AOI22_X1 U1086 ( .A1(\REGISTERS[28][18] ), .A2(n108), .B1(
        \REGISTERS[29][18] ), .B2(n1489), .ZN(n1043) );
  AOI22_X1 U1087 ( .A1(\REGISTERS[30][18] ), .A2(n110), .B1(\REGISTERS[7][18] ), .B2(n1491), .ZN(n1042) );
  AOI22_X1 U1088 ( .A1(\REGISTERS[5][18] ), .A2(n112), .B1(\REGISTERS[3][18] ), 
        .B2(n1493), .ZN(n1041) );
  NAND4_X1 U1089 ( .A1(n1044), .A2(n1043), .A3(n1042), .A4(n1041), .ZN(n1056)
         );
  AOI22_X1 U1090 ( .A1(\REGISTERS[9][18] ), .A2(n114), .B1(\REGISTERS[10][18] ), .B2(n113), .ZN(n1048) );
  AOI22_X1 U1091 ( .A1(\REGISTERS[11][18] ), .A2(n116), .B1(
        \REGISTERS[12][18] ), .B2(n115), .ZN(n1047) );
  AOI22_X1 U1092 ( .A1(\REGISTERS[13][18] ), .A2(n118), .B1(
        \REGISTERS[14][18] ), .B2(n117), .ZN(n1046) );
  AOI22_X1 U1093 ( .A1(\REGISTERS[15][18] ), .A2(n120), .B1(
        \REGISTERS[17][18] ), .B2(n119), .ZN(n1045) );
  NAND4_X1 U1094 ( .A1(n1048), .A2(n1047), .A3(n1046), .A4(n1045), .ZN(n1055)
         );
  AOI22_X1 U1095 ( .A1(\REGISTERS[31][18] ), .A2(n122), .B1(
        \REGISTERS[22][18] ), .B2(n1511), .ZN(n1049) );
  OAI21_X1 U1096 ( .B1(n47), .B2(n1514), .A(n1049), .ZN(n1054) );
  AOI22_X1 U1097 ( .A1(\REGISTERS[24][18] ), .A2(n124), .B1(
        \REGISTERS[25][18] ), .B2(n1515), .ZN(n1052) );
  AOI22_X1 U1098 ( .A1(\REGISTERS[8][18] ), .A2(n36), .B1(\REGISTERS[23][18] ), 
        .B2(n125), .ZN(n1051) );
  AOI22_X1 U1099 ( .A1(\REGISTERS[16][18] ), .A2(n1520), .B1(
        \REGISTERS[1][18] ), .B2(n37), .ZN(n1050) );
  NAND3_X1 U1100 ( .A1(n1052), .A2(n1051), .A3(n1050), .ZN(n1053) );
  NOR4_X1 U1101 ( .A1(n1056), .A2(n1055), .A3(n1054), .A4(n1053), .ZN(n1057)
         );
  NAND4_X1 U1102 ( .A1(n1060), .A2(n1059), .A3(n1058), .A4(n1057), .ZN(
        OUT2[18]) );
  AOI22_X1 U1103 ( .A1(\REGISTERS[18][19] ), .A2(n100), .B1(
        \REGISTERS[19][19] ), .B2(n1481), .ZN(n1080) );
  AOI22_X1 U1104 ( .A1(\REGISTERS[20][19] ), .A2(n102), .B1(
        \REGISTERS[21][19] ), .B2(n1483), .ZN(n1079) );
  AOI22_X1 U1105 ( .A1(\REGISTERS[4][19] ), .A2(n104), .B1(\REGISTERS[2][19] ), 
        .B2(n1485), .ZN(n1078) );
  AOI22_X1 U1106 ( .A1(\REGISTERS[26][19] ), .A2(n106), .B1(
        \REGISTERS[27][19] ), .B2(n1487), .ZN(n1064) );
  AOI22_X1 U1107 ( .A1(\REGISTERS[28][19] ), .A2(n108), .B1(
        \REGISTERS[29][19] ), .B2(n1489), .ZN(n1063) );
  AOI22_X1 U1108 ( .A1(\REGISTERS[30][19] ), .A2(n110), .B1(\REGISTERS[7][19] ), .B2(n1491), .ZN(n1062) );
  AOI22_X1 U1109 ( .A1(\REGISTERS[5][19] ), .A2(n112), .B1(\REGISTERS[3][19] ), 
        .B2(n1493), .ZN(n1061) );
  NAND4_X1 U1110 ( .A1(n1064), .A2(n1063), .A3(n1062), .A4(n1061), .ZN(n1076)
         );
  AOI22_X1 U1111 ( .A1(\REGISTERS[9][19] ), .A2(n114), .B1(\REGISTERS[10][19] ), .B2(n1499), .ZN(n1068) );
  AOI22_X1 U1112 ( .A1(\REGISTERS[11][19] ), .A2(n116), .B1(
        \REGISTERS[12][19] ), .B2(n1501), .ZN(n1067) );
  AOI22_X1 U1113 ( .A1(\REGISTERS[13][19] ), .A2(n118), .B1(
        \REGISTERS[14][19] ), .B2(n1503), .ZN(n1066) );
  AOI22_X1 U1114 ( .A1(\REGISTERS[15][19] ), .A2(n120), .B1(
        \REGISTERS[17][19] ), .B2(n1505), .ZN(n1065) );
  NAND4_X1 U1115 ( .A1(n1068), .A2(n1067), .A3(n1066), .A4(n1065), .ZN(n1075)
         );
  AOI22_X1 U1116 ( .A1(\REGISTERS[31][19] ), .A2(n122), .B1(
        \REGISTERS[22][19] ), .B2(n121), .ZN(n1069) );
  OAI21_X1 U1117 ( .B1(n48), .B2(n1514), .A(n1069), .ZN(n1074) );
  AOI22_X1 U1118 ( .A1(\REGISTERS[24][19] ), .A2(n124), .B1(
        \REGISTERS[25][19] ), .B2(n1515), .ZN(n1072) );
  AOI22_X1 U1119 ( .A1(\REGISTERS[8][19] ), .A2(n36), .B1(\REGISTERS[23][19] ), 
        .B2(n1517), .ZN(n1071) );
  AOI22_X1 U1120 ( .A1(\REGISTERS[16][19] ), .A2(n1520), .B1(
        \REGISTERS[1][19] ), .B2(n37), .ZN(n1070) );
  NAND3_X1 U1121 ( .A1(n1072), .A2(n1071), .A3(n1070), .ZN(n1073) );
  NOR4_X1 U1122 ( .A1(n1076), .A2(n1075), .A3(n1074), .A4(n1073), .ZN(n1077)
         );
  NAND4_X1 U1123 ( .A1(n1080), .A2(n1079), .A3(n1078), .A4(n1077), .ZN(
        OUT2[19]) );
  AOI22_X1 U1124 ( .A1(\REGISTERS[18][1] ), .A2(n100), .B1(\REGISTERS[19][1] ), 
        .B2(n99), .ZN(n1100) );
  AOI22_X1 U1125 ( .A1(\REGISTERS[20][1] ), .A2(n102), .B1(\REGISTERS[21][1] ), 
        .B2(n101), .ZN(n1099) );
  AOI22_X1 U1126 ( .A1(\REGISTERS[4][1] ), .A2(n104), .B1(\REGISTERS[2][1] ), 
        .B2(n103), .ZN(n1098) );
  AOI22_X1 U1127 ( .A1(\REGISTERS[26][1] ), .A2(n106), .B1(\REGISTERS[27][1] ), 
        .B2(n105), .ZN(n1084) );
  AOI22_X1 U1128 ( .A1(\REGISTERS[28][1] ), .A2(n108), .B1(\REGISTERS[29][1] ), 
        .B2(n107), .ZN(n1083) );
  AOI22_X1 U1129 ( .A1(\REGISTERS[30][1] ), .A2(n110), .B1(\REGISTERS[7][1] ), 
        .B2(n109), .ZN(n1082) );
  AOI22_X1 U1130 ( .A1(\REGISTERS[5][1] ), .A2(n112), .B1(\REGISTERS[3][1] ), 
        .B2(n111), .ZN(n1081) );
  NAND4_X1 U1131 ( .A1(n1084), .A2(n1083), .A3(n1082), .A4(n1081), .ZN(n1096)
         );
  AOI22_X1 U1132 ( .A1(\REGISTERS[9][1] ), .A2(n114), .B1(\REGISTERS[10][1] ), 
        .B2(n113), .ZN(n1088) );
  AOI22_X1 U1133 ( .A1(\REGISTERS[11][1] ), .A2(n116), .B1(\REGISTERS[12][1] ), 
        .B2(n115), .ZN(n1087) );
  AOI22_X1 U1134 ( .A1(\REGISTERS[13][1] ), .A2(n118), .B1(\REGISTERS[14][1] ), 
        .B2(n117), .ZN(n1086) );
  AOI22_X1 U1135 ( .A1(\REGISTERS[15][1] ), .A2(n120), .B1(\REGISTERS[17][1] ), 
        .B2(n119), .ZN(n1085) );
  NAND4_X1 U1136 ( .A1(n1088), .A2(n1087), .A3(n1086), .A4(n1085), .ZN(n1095)
         );
  AOI22_X1 U1137 ( .A1(\REGISTERS[31][1] ), .A2(n122), .B1(\REGISTERS[22][1] ), 
        .B2(n121), .ZN(n1089) );
  OAI21_X1 U1138 ( .B1(n49), .B2(n1514), .A(n1089), .ZN(n1094) );
  AOI22_X1 U1139 ( .A1(\REGISTERS[24][1] ), .A2(n124), .B1(\REGISTERS[25][1] ), 
        .B2(n123), .ZN(n1092) );
  AOI22_X1 U1140 ( .A1(\REGISTERS[8][1] ), .A2(n36), .B1(\REGISTERS[23][1] ), 
        .B2(n125), .ZN(n1091) );
  AOI22_X1 U1141 ( .A1(\REGISTERS[16][1] ), .A2(n1520), .B1(\REGISTERS[1][1] ), 
        .B2(n37), .ZN(n1090) );
  NAND3_X1 U1142 ( .A1(n1092), .A2(n1091), .A3(n1090), .ZN(n1093) );
  NOR4_X1 U1143 ( .A1(n1096), .A2(n1095), .A3(n1094), .A4(n1093), .ZN(n1097)
         );
  NAND4_X1 U1144 ( .A1(n1100), .A2(n1099), .A3(n1098), .A4(n1097), .ZN(OUT2[1]) );
  AOI22_X1 U1145 ( .A1(\REGISTERS[18][20] ), .A2(n100), .B1(
        \REGISTERS[19][20] ), .B2(n99), .ZN(n1120) );
  AOI22_X1 U1146 ( .A1(\REGISTERS[20][20] ), .A2(n102), .B1(
        \REGISTERS[21][20] ), .B2(n101), .ZN(n1119) );
  AOI22_X1 U1147 ( .A1(\REGISTERS[4][20] ), .A2(n104), .B1(\REGISTERS[2][20] ), 
        .B2(n103), .ZN(n1118) );
  AOI22_X1 U1148 ( .A1(\REGISTERS[26][20] ), .A2(n106), .B1(
        \REGISTERS[27][20] ), .B2(n105), .ZN(n1104) );
  AOI22_X1 U1149 ( .A1(\REGISTERS[28][20] ), .A2(n108), .B1(
        \REGISTERS[29][20] ), .B2(n107), .ZN(n1103) );
  AOI22_X1 U1150 ( .A1(\REGISTERS[30][20] ), .A2(n110), .B1(\REGISTERS[7][20] ), .B2(n109), .ZN(n1102) );
  AOI22_X1 U1151 ( .A1(\REGISTERS[5][20] ), .A2(n112), .B1(\REGISTERS[3][20] ), 
        .B2(n111), .ZN(n1101) );
  NAND4_X1 U1152 ( .A1(n1104), .A2(n1103), .A3(n1102), .A4(n1101), .ZN(n1116)
         );
  AOI22_X1 U1153 ( .A1(\REGISTERS[9][20] ), .A2(n114), .B1(\REGISTERS[10][20] ), .B2(n113), .ZN(n1108) );
  AOI22_X1 U1154 ( .A1(\REGISTERS[11][20] ), .A2(n116), .B1(
        \REGISTERS[12][20] ), .B2(n115), .ZN(n1107) );
  AOI22_X1 U1155 ( .A1(\REGISTERS[13][20] ), .A2(n118), .B1(
        \REGISTERS[14][20] ), .B2(n117), .ZN(n1106) );
  AOI22_X1 U1156 ( .A1(\REGISTERS[15][20] ), .A2(n120), .B1(
        \REGISTERS[17][20] ), .B2(n119), .ZN(n1105) );
  NAND4_X1 U1157 ( .A1(n1108), .A2(n1107), .A3(n1106), .A4(n1105), .ZN(n1115)
         );
  AOI22_X1 U1158 ( .A1(\REGISTERS[31][20] ), .A2(n122), .B1(
        \REGISTERS[22][20] ), .B2(n121), .ZN(n1109) );
  OAI21_X1 U1159 ( .B1(n50), .B2(n1514), .A(n1109), .ZN(n1114) );
  AOI22_X1 U1160 ( .A1(\REGISTERS[24][20] ), .A2(n124), .B1(
        \REGISTERS[25][20] ), .B2(n123), .ZN(n1112) );
  AOI22_X1 U1161 ( .A1(\REGISTERS[8][20] ), .A2(n36), .B1(\REGISTERS[23][20] ), 
        .B2(n125), .ZN(n1111) );
  AOI22_X1 U1162 ( .A1(\REGISTERS[16][20] ), .A2(n1520), .B1(
        \REGISTERS[1][20] ), .B2(n37), .ZN(n1110) );
  NAND3_X1 U1163 ( .A1(n1112), .A2(n1111), .A3(n1110), .ZN(n1113) );
  NOR4_X1 U1164 ( .A1(n1116), .A2(n1115), .A3(n1114), .A4(n1113), .ZN(n1117)
         );
  NAND4_X1 U1165 ( .A1(n1120), .A2(n1119), .A3(n1118), .A4(n1117), .ZN(
        OUT2[20]) );
  AOI22_X1 U1166 ( .A1(\REGISTERS[18][21] ), .A2(n100), .B1(
        \REGISTERS[19][21] ), .B2(n99), .ZN(n1140) );
  AOI22_X1 U1167 ( .A1(\REGISTERS[20][21] ), .A2(n102), .B1(
        \REGISTERS[21][21] ), .B2(n101), .ZN(n1139) );
  AOI22_X1 U1168 ( .A1(\REGISTERS[4][21] ), .A2(n104), .B1(\REGISTERS[2][21] ), 
        .B2(n103), .ZN(n1138) );
  AOI22_X1 U1169 ( .A1(\REGISTERS[26][21] ), .A2(n106), .B1(
        \REGISTERS[27][21] ), .B2(n105), .ZN(n1124) );
  AOI22_X1 U1170 ( .A1(\REGISTERS[28][21] ), .A2(n108), .B1(
        \REGISTERS[29][21] ), .B2(n107), .ZN(n1123) );
  AOI22_X1 U1171 ( .A1(\REGISTERS[30][21] ), .A2(n110), .B1(\REGISTERS[7][21] ), .B2(n109), .ZN(n1122) );
  AOI22_X1 U1172 ( .A1(\REGISTERS[5][21] ), .A2(n112), .B1(\REGISTERS[3][21] ), 
        .B2(n111), .ZN(n1121) );
  NAND4_X1 U1173 ( .A1(n1124), .A2(n1123), .A3(n1122), .A4(n1121), .ZN(n1136)
         );
  AOI22_X1 U1174 ( .A1(\REGISTERS[9][21] ), .A2(n114), .B1(\REGISTERS[10][21] ), .B2(n113), .ZN(n1128) );
  AOI22_X1 U1175 ( .A1(\REGISTERS[11][21] ), .A2(n116), .B1(
        \REGISTERS[12][21] ), .B2(n115), .ZN(n1127) );
  AOI22_X1 U1176 ( .A1(\REGISTERS[13][21] ), .A2(n118), .B1(
        \REGISTERS[14][21] ), .B2(n117), .ZN(n1126) );
  AOI22_X1 U1177 ( .A1(\REGISTERS[15][21] ), .A2(n120), .B1(
        \REGISTERS[17][21] ), .B2(n119), .ZN(n1125) );
  NAND4_X1 U1178 ( .A1(n1128), .A2(n1127), .A3(n1126), .A4(n1125), .ZN(n1135)
         );
  AOI22_X1 U1179 ( .A1(\REGISTERS[31][21] ), .A2(n122), .B1(
        \REGISTERS[22][21] ), .B2(n121), .ZN(n1129) );
  OAI21_X1 U1180 ( .B1(n51), .B2(n1514), .A(n1129), .ZN(n1134) );
  AOI22_X1 U1181 ( .A1(\REGISTERS[24][21] ), .A2(n124), .B1(
        \REGISTERS[25][21] ), .B2(n123), .ZN(n1132) );
  AOI22_X1 U1182 ( .A1(\REGISTERS[8][21] ), .A2(n36), .B1(\REGISTERS[23][21] ), 
        .B2(n125), .ZN(n1131) );
  AOI22_X1 U1183 ( .A1(\REGISTERS[16][21] ), .A2(n1520), .B1(
        \REGISTERS[1][21] ), .B2(n37), .ZN(n1130) );
  NAND3_X1 U1184 ( .A1(n1132), .A2(n1131), .A3(n1130), .ZN(n1133) );
  NOR4_X1 U1185 ( .A1(n1136), .A2(n1135), .A3(n1134), .A4(n1133), .ZN(n1137)
         );
  NAND4_X1 U1186 ( .A1(n1140), .A2(n1139), .A3(n1138), .A4(n1137), .ZN(
        OUT2[21]) );
  AOI22_X1 U1187 ( .A1(\REGISTERS[18][22] ), .A2(n100), .B1(
        \REGISTERS[19][22] ), .B2(n99), .ZN(n1160) );
  AOI22_X1 U1188 ( .A1(\REGISTERS[20][22] ), .A2(n102), .B1(
        \REGISTERS[21][22] ), .B2(n101), .ZN(n1159) );
  AOI22_X1 U1189 ( .A1(\REGISTERS[4][22] ), .A2(n104), .B1(\REGISTERS[2][22] ), 
        .B2(n103), .ZN(n1158) );
  AOI22_X1 U1190 ( .A1(\REGISTERS[26][22] ), .A2(n106), .B1(
        \REGISTERS[27][22] ), .B2(n105), .ZN(n1144) );
  AOI22_X1 U1191 ( .A1(\REGISTERS[28][22] ), .A2(n108), .B1(
        \REGISTERS[29][22] ), .B2(n107), .ZN(n1143) );
  AOI22_X1 U1192 ( .A1(\REGISTERS[30][22] ), .A2(n110), .B1(\REGISTERS[7][22] ), .B2(n109), .ZN(n1142) );
  AOI22_X1 U1193 ( .A1(\REGISTERS[5][22] ), .A2(n112), .B1(\REGISTERS[3][22] ), 
        .B2(n111), .ZN(n1141) );
  NAND4_X1 U1194 ( .A1(n1144), .A2(n1143), .A3(n1142), .A4(n1141), .ZN(n1156)
         );
  AOI22_X1 U1195 ( .A1(\REGISTERS[9][22] ), .A2(n114), .B1(\REGISTERS[10][22] ), .B2(n113), .ZN(n1148) );
  AOI22_X1 U1196 ( .A1(\REGISTERS[11][22] ), .A2(n116), .B1(
        \REGISTERS[12][22] ), .B2(n115), .ZN(n1147) );
  AOI22_X1 U1197 ( .A1(\REGISTERS[13][22] ), .A2(n118), .B1(
        \REGISTERS[14][22] ), .B2(n117), .ZN(n1146) );
  AOI22_X1 U1198 ( .A1(\REGISTERS[15][22] ), .A2(n120), .B1(
        \REGISTERS[17][22] ), .B2(n119), .ZN(n1145) );
  NAND4_X1 U1199 ( .A1(n1148), .A2(n1147), .A3(n1146), .A4(n1145), .ZN(n1155)
         );
  AOI22_X1 U1200 ( .A1(\REGISTERS[31][22] ), .A2(n122), .B1(
        \REGISTERS[22][22] ), .B2(n121), .ZN(n1149) );
  OAI21_X1 U1201 ( .B1(n52), .B2(n1514), .A(n1149), .ZN(n1154) );
  AOI22_X1 U1202 ( .A1(\REGISTERS[24][22] ), .A2(n124), .B1(
        \REGISTERS[25][22] ), .B2(n123), .ZN(n1152) );
  AOI22_X1 U1203 ( .A1(\REGISTERS[8][22] ), .A2(n36), .B1(\REGISTERS[23][22] ), 
        .B2(n125), .ZN(n1151) );
  AOI22_X1 U1204 ( .A1(\REGISTERS[16][22] ), .A2(n1520), .B1(
        \REGISTERS[1][22] ), .B2(n37), .ZN(n1150) );
  NAND3_X1 U1205 ( .A1(n1152), .A2(n1151), .A3(n1150), .ZN(n1153) );
  NOR4_X1 U1206 ( .A1(n1156), .A2(n1155), .A3(n1154), .A4(n1153), .ZN(n1157)
         );
  NAND4_X1 U1207 ( .A1(n1160), .A2(n1159), .A3(n1158), .A4(n1157), .ZN(
        OUT2[22]) );
  AOI22_X1 U1208 ( .A1(\REGISTERS[18][23] ), .A2(n100), .B1(
        \REGISTERS[19][23] ), .B2(n99), .ZN(n1180) );
  AOI22_X1 U1209 ( .A1(\REGISTERS[20][23] ), .A2(n102), .B1(
        \REGISTERS[21][23] ), .B2(n101), .ZN(n1179) );
  AOI22_X1 U1210 ( .A1(\REGISTERS[4][23] ), .A2(n104), .B1(\REGISTERS[2][23] ), 
        .B2(n103), .ZN(n1178) );
  AOI22_X1 U1211 ( .A1(\REGISTERS[26][23] ), .A2(n106), .B1(
        \REGISTERS[27][23] ), .B2(n105), .ZN(n1164) );
  AOI22_X1 U1212 ( .A1(\REGISTERS[28][23] ), .A2(n108), .B1(
        \REGISTERS[29][23] ), .B2(n107), .ZN(n1163) );
  AOI22_X1 U1213 ( .A1(\REGISTERS[30][23] ), .A2(n110), .B1(\REGISTERS[7][23] ), .B2(n109), .ZN(n1162) );
  AOI22_X1 U1214 ( .A1(\REGISTERS[5][23] ), .A2(n112), .B1(\REGISTERS[3][23] ), 
        .B2(n111), .ZN(n1161) );
  NAND4_X1 U1215 ( .A1(n1164), .A2(n1163), .A3(n1162), .A4(n1161), .ZN(n1176)
         );
  AOI22_X1 U1216 ( .A1(\REGISTERS[9][23] ), .A2(n114), .B1(\REGISTERS[10][23] ), .B2(n113), .ZN(n1168) );
  AOI22_X1 U1217 ( .A1(\REGISTERS[11][23] ), .A2(n116), .B1(
        \REGISTERS[12][23] ), .B2(n115), .ZN(n1167) );
  AOI22_X1 U1218 ( .A1(\REGISTERS[13][23] ), .A2(n118), .B1(
        \REGISTERS[14][23] ), .B2(n117), .ZN(n1166) );
  AOI22_X1 U1219 ( .A1(\REGISTERS[15][23] ), .A2(n120), .B1(
        \REGISTERS[17][23] ), .B2(n119), .ZN(n1165) );
  NAND4_X1 U1220 ( .A1(n1168), .A2(n1167), .A3(n1166), .A4(n1165), .ZN(n1175)
         );
  AOI22_X1 U1221 ( .A1(\REGISTERS[31][23] ), .A2(n122), .B1(
        \REGISTERS[22][23] ), .B2(n121), .ZN(n1169) );
  OAI21_X1 U1222 ( .B1(n53), .B2(n1514), .A(n1169), .ZN(n1174) );
  AOI22_X1 U1223 ( .A1(\REGISTERS[24][23] ), .A2(n124), .B1(
        \REGISTERS[25][23] ), .B2(n123), .ZN(n1172) );
  AOI22_X1 U1224 ( .A1(\REGISTERS[8][23] ), .A2(n36), .B1(\REGISTERS[23][23] ), 
        .B2(n125), .ZN(n1171) );
  AOI22_X1 U1225 ( .A1(\REGISTERS[16][23] ), .A2(n1520), .B1(
        \REGISTERS[1][23] ), .B2(n37), .ZN(n1170) );
  NAND3_X1 U1226 ( .A1(n1172), .A2(n1171), .A3(n1170), .ZN(n1173) );
  NOR4_X1 U1227 ( .A1(n1176), .A2(n1175), .A3(n1174), .A4(n1173), .ZN(n1177)
         );
  NAND4_X1 U1228 ( .A1(n1180), .A2(n1179), .A3(n1178), .A4(n1177), .ZN(
        OUT2[23]) );
  AOI22_X1 U1229 ( .A1(\REGISTERS[18][24] ), .A2(n100), .B1(
        \REGISTERS[19][24] ), .B2(n99), .ZN(n1200) );
  AOI22_X1 U1230 ( .A1(\REGISTERS[20][24] ), .A2(n102), .B1(
        \REGISTERS[21][24] ), .B2(n101), .ZN(n1199) );
  AOI22_X1 U1231 ( .A1(\REGISTERS[4][24] ), .A2(n104), .B1(\REGISTERS[2][24] ), 
        .B2(n103), .ZN(n1198) );
  AOI22_X1 U1232 ( .A1(\REGISTERS[26][24] ), .A2(n106), .B1(
        \REGISTERS[27][24] ), .B2(n105), .ZN(n1184) );
  AOI22_X1 U1233 ( .A1(\REGISTERS[28][24] ), .A2(n108), .B1(
        \REGISTERS[29][24] ), .B2(n107), .ZN(n1183) );
  AOI22_X1 U1234 ( .A1(\REGISTERS[30][24] ), .A2(n110), .B1(\REGISTERS[7][24] ), .B2(n109), .ZN(n1182) );
  AOI22_X1 U1235 ( .A1(\REGISTERS[5][24] ), .A2(n112), .B1(\REGISTERS[3][24] ), 
        .B2(n111), .ZN(n1181) );
  NAND4_X1 U1236 ( .A1(n1184), .A2(n1183), .A3(n1182), .A4(n1181), .ZN(n1196)
         );
  AOI22_X1 U1237 ( .A1(\REGISTERS[9][24] ), .A2(n114), .B1(\REGISTERS[10][24] ), .B2(n113), .ZN(n1188) );
  AOI22_X1 U1238 ( .A1(\REGISTERS[11][24] ), .A2(n116), .B1(
        \REGISTERS[12][24] ), .B2(n115), .ZN(n1187) );
  AOI22_X1 U1239 ( .A1(\REGISTERS[13][24] ), .A2(n118), .B1(
        \REGISTERS[14][24] ), .B2(n117), .ZN(n1186) );
  AOI22_X1 U1240 ( .A1(\REGISTERS[15][24] ), .A2(n120), .B1(
        \REGISTERS[17][24] ), .B2(n119), .ZN(n1185) );
  NAND4_X1 U1241 ( .A1(n1188), .A2(n1187), .A3(n1186), .A4(n1185), .ZN(n1195)
         );
  AOI22_X1 U1242 ( .A1(\REGISTERS[31][24] ), .A2(n122), .B1(
        \REGISTERS[22][24] ), .B2(n121), .ZN(n1189) );
  OAI21_X1 U1243 ( .B1(n54), .B2(n1514), .A(n1189), .ZN(n1194) );
  AOI22_X1 U1244 ( .A1(\REGISTERS[24][24] ), .A2(n124), .B1(
        \REGISTERS[25][24] ), .B2(n123), .ZN(n1192) );
  AOI22_X1 U1245 ( .A1(\REGISTERS[8][24] ), .A2(n36), .B1(\REGISTERS[23][24] ), 
        .B2(n125), .ZN(n1191) );
  AOI22_X1 U1246 ( .A1(\REGISTERS[16][24] ), .A2(n1520), .B1(
        \REGISTERS[1][24] ), .B2(n37), .ZN(n1190) );
  NAND3_X1 U1247 ( .A1(n1192), .A2(n1191), .A3(n1190), .ZN(n1193) );
  NOR4_X1 U1248 ( .A1(n1196), .A2(n1195), .A3(n1194), .A4(n1193), .ZN(n1197)
         );
  NAND4_X1 U1249 ( .A1(n1200), .A2(n1199), .A3(n1198), .A4(n1197), .ZN(
        OUT2[24]) );
  AOI22_X1 U1250 ( .A1(\REGISTERS[18][25] ), .A2(n100), .B1(
        \REGISTERS[19][25] ), .B2(n99), .ZN(n1220) );
  AOI22_X1 U1251 ( .A1(\REGISTERS[20][25] ), .A2(n102), .B1(
        \REGISTERS[21][25] ), .B2(n101), .ZN(n1219) );
  AOI22_X1 U1252 ( .A1(\REGISTERS[4][25] ), .A2(n104), .B1(\REGISTERS[2][25] ), 
        .B2(n103), .ZN(n1218) );
  AOI22_X1 U1253 ( .A1(\REGISTERS[26][25] ), .A2(n106), .B1(
        \REGISTERS[27][25] ), .B2(n105), .ZN(n1204) );
  AOI22_X1 U1254 ( .A1(\REGISTERS[28][25] ), .A2(n108), .B1(
        \REGISTERS[29][25] ), .B2(n107), .ZN(n1203) );
  AOI22_X1 U1255 ( .A1(\REGISTERS[30][25] ), .A2(n110), .B1(\REGISTERS[7][25] ), .B2(n109), .ZN(n1202) );
  AOI22_X1 U1256 ( .A1(\REGISTERS[5][25] ), .A2(n112), .B1(\REGISTERS[3][25] ), 
        .B2(n111), .ZN(n1201) );
  NAND4_X1 U1257 ( .A1(n1204), .A2(n1203), .A3(n1202), .A4(n1201), .ZN(n1216)
         );
  AOI22_X1 U1258 ( .A1(\REGISTERS[9][25] ), .A2(n114), .B1(\REGISTERS[10][25] ), .B2(n113), .ZN(n1208) );
  AOI22_X1 U1259 ( .A1(\REGISTERS[11][25] ), .A2(n116), .B1(
        \REGISTERS[12][25] ), .B2(n115), .ZN(n1207) );
  AOI22_X1 U1260 ( .A1(\REGISTERS[13][25] ), .A2(n118), .B1(
        \REGISTERS[14][25] ), .B2(n117), .ZN(n1206) );
  AOI22_X1 U1261 ( .A1(\REGISTERS[15][25] ), .A2(n120), .B1(
        \REGISTERS[17][25] ), .B2(n119), .ZN(n1205) );
  NAND4_X1 U1262 ( .A1(n1208), .A2(n1207), .A3(n1206), .A4(n1205), .ZN(n1215)
         );
  AOI22_X1 U1263 ( .A1(\REGISTERS[31][25] ), .A2(n122), .B1(
        \REGISTERS[22][25] ), .B2(n121), .ZN(n1209) );
  OAI21_X1 U1264 ( .B1(n55), .B2(n1514), .A(n1209), .ZN(n1214) );
  AOI22_X1 U1265 ( .A1(\REGISTERS[24][25] ), .A2(n124), .B1(
        \REGISTERS[25][25] ), .B2(n123), .ZN(n1212) );
  AOI22_X1 U1266 ( .A1(\REGISTERS[8][25] ), .A2(n36), .B1(\REGISTERS[23][25] ), 
        .B2(n125), .ZN(n1211) );
  AOI22_X1 U1267 ( .A1(\REGISTERS[16][25] ), .A2(n1520), .B1(
        \REGISTERS[1][25] ), .B2(n37), .ZN(n1210) );
  NAND3_X1 U1268 ( .A1(n1212), .A2(n1211), .A3(n1210), .ZN(n1213) );
  NOR4_X1 U1269 ( .A1(n1216), .A2(n1215), .A3(n1214), .A4(n1213), .ZN(n1217)
         );
  NAND4_X1 U1270 ( .A1(n1220), .A2(n1219), .A3(n1218), .A4(n1217), .ZN(
        OUT2[25]) );
  AOI22_X1 U1271 ( .A1(\REGISTERS[18][26] ), .A2(n100), .B1(
        \REGISTERS[19][26] ), .B2(n99), .ZN(n1240) );
  AOI22_X1 U1272 ( .A1(\REGISTERS[20][26] ), .A2(n102), .B1(
        \REGISTERS[21][26] ), .B2(n101), .ZN(n1239) );
  AOI22_X1 U1273 ( .A1(\REGISTERS[4][26] ), .A2(n104), .B1(\REGISTERS[2][26] ), 
        .B2(n103), .ZN(n1238) );
  AOI22_X1 U1274 ( .A1(\REGISTERS[26][26] ), .A2(n106), .B1(
        \REGISTERS[27][26] ), .B2(n105), .ZN(n1224) );
  AOI22_X1 U1275 ( .A1(\REGISTERS[28][26] ), .A2(n108), .B1(
        \REGISTERS[29][26] ), .B2(n107), .ZN(n1223) );
  AOI22_X1 U1276 ( .A1(\REGISTERS[30][26] ), .A2(n110), .B1(\REGISTERS[7][26] ), .B2(n109), .ZN(n1222) );
  AOI22_X1 U1277 ( .A1(\REGISTERS[5][26] ), .A2(n112), .B1(\REGISTERS[3][26] ), 
        .B2(n111), .ZN(n1221) );
  NAND4_X1 U1278 ( .A1(n1224), .A2(n1223), .A3(n1222), .A4(n1221), .ZN(n1236)
         );
  AOI22_X1 U1279 ( .A1(\REGISTERS[9][26] ), .A2(n114), .B1(\REGISTERS[10][26] ), .B2(n113), .ZN(n1228) );
  AOI22_X1 U1280 ( .A1(\REGISTERS[11][26] ), .A2(n116), .B1(
        \REGISTERS[12][26] ), .B2(n115), .ZN(n1227) );
  AOI22_X1 U1281 ( .A1(\REGISTERS[13][26] ), .A2(n118), .B1(
        \REGISTERS[14][26] ), .B2(n117), .ZN(n1226) );
  AOI22_X1 U1282 ( .A1(\REGISTERS[15][26] ), .A2(n120), .B1(
        \REGISTERS[17][26] ), .B2(n119), .ZN(n1225) );
  NAND4_X1 U1283 ( .A1(n1228), .A2(n1227), .A3(n1226), .A4(n1225), .ZN(n1235)
         );
  AOI22_X1 U1284 ( .A1(\REGISTERS[31][26] ), .A2(n122), .B1(
        \REGISTERS[22][26] ), .B2(n121), .ZN(n1229) );
  OAI21_X1 U1285 ( .B1(n56), .B2(n1514), .A(n1229), .ZN(n1234) );
  AOI22_X1 U1286 ( .A1(\REGISTERS[24][26] ), .A2(n124), .B1(
        \REGISTERS[25][26] ), .B2(n123), .ZN(n1232) );
  AOI22_X1 U1287 ( .A1(\REGISTERS[8][26] ), .A2(n36), .B1(\REGISTERS[23][26] ), 
        .B2(n125), .ZN(n1231) );
  AOI22_X1 U1288 ( .A1(\REGISTERS[16][26] ), .A2(n1520), .B1(
        \REGISTERS[1][26] ), .B2(n37), .ZN(n1230) );
  NAND3_X1 U1289 ( .A1(n1232), .A2(n1231), .A3(n1230), .ZN(n1233) );
  NOR4_X1 U1290 ( .A1(n1236), .A2(n1235), .A3(n1234), .A4(n1233), .ZN(n1237)
         );
  NAND4_X1 U1291 ( .A1(n1240), .A2(n1239), .A3(n1238), .A4(n1237), .ZN(
        OUT2[26]) );
  AOI22_X1 U1292 ( .A1(\REGISTERS[18][27] ), .A2(n100), .B1(
        \REGISTERS[19][27] ), .B2(n99), .ZN(n1260) );
  AOI22_X1 U1293 ( .A1(\REGISTERS[20][27] ), .A2(n102), .B1(
        \REGISTERS[21][27] ), .B2(n101), .ZN(n1259) );
  AOI22_X1 U1294 ( .A1(\REGISTERS[4][27] ), .A2(n104), .B1(\REGISTERS[2][27] ), 
        .B2(n103), .ZN(n1258) );
  AOI22_X1 U1295 ( .A1(\REGISTERS[26][27] ), .A2(n106), .B1(
        \REGISTERS[27][27] ), .B2(n105), .ZN(n1244) );
  AOI22_X1 U1296 ( .A1(\REGISTERS[28][27] ), .A2(n108), .B1(
        \REGISTERS[29][27] ), .B2(n107), .ZN(n1243) );
  AOI22_X1 U1297 ( .A1(\REGISTERS[30][27] ), .A2(n110), .B1(\REGISTERS[7][27] ), .B2(n109), .ZN(n1242) );
  AOI22_X1 U1298 ( .A1(\REGISTERS[5][27] ), .A2(n1494), .B1(\REGISTERS[3][27] ), .B2(n111), .ZN(n1241) );
  NAND4_X1 U1299 ( .A1(n1244), .A2(n1243), .A3(n1242), .A4(n1241), .ZN(n1256)
         );
  AOI22_X1 U1300 ( .A1(\REGISTERS[9][27] ), .A2(n114), .B1(\REGISTERS[10][27] ), .B2(n113), .ZN(n1248) );
  AOI22_X1 U1301 ( .A1(\REGISTERS[11][27] ), .A2(n116), .B1(
        \REGISTERS[12][27] ), .B2(n115), .ZN(n1247) );
  AOI22_X1 U1302 ( .A1(\REGISTERS[13][27] ), .A2(n118), .B1(
        \REGISTERS[14][27] ), .B2(n117), .ZN(n1246) );
  AOI22_X1 U1303 ( .A1(\REGISTERS[15][27] ), .A2(n120), .B1(
        \REGISTERS[17][27] ), .B2(n119), .ZN(n1245) );
  NAND4_X1 U1304 ( .A1(n1248), .A2(n1247), .A3(n1246), .A4(n1245), .ZN(n1255)
         );
  AOI22_X1 U1305 ( .A1(\REGISTERS[31][27] ), .A2(n122), .B1(
        \REGISTERS[22][27] ), .B2(n121), .ZN(n1249) );
  OAI21_X1 U1306 ( .B1(n57), .B2(n1514), .A(n1249), .ZN(n1254) );
  AOI22_X1 U1307 ( .A1(\REGISTERS[24][27] ), .A2(n124), .B1(
        \REGISTERS[25][27] ), .B2(n123), .ZN(n1252) );
  AOI22_X1 U1308 ( .A1(\REGISTERS[8][27] ), .A2(n36), .B1(\REGISTERS[23][27] ), 
        .B2(n125), .ZN(n1251) );
  AOI22_X1 U1309 ( .A1(\REGISTERS[16][27] ), .A2(n1520), .B1(
        \REGISTERS[1][27] ), .B2(n37), .ZN(n1250) );
  NAND3_X1 U1310 ( .A1(n1252), .A2(n1251), .A3(n1250), .ZN(n1253) );
  NOR4_X1 U1311 ( .A1(n1256), .A2(n1255), .A3(n1254), .A4(n1253), .ZN(n1257)
         );
  NAND4_X1 U1312 ( .A1(n1260), .A2(n1259), .A3(n1258), .A4(n1257), .ZN(
        OUT2[27]) );
  AOI22_X1 U1313 ( .A1(\REGISTERS[18][28] ), .A2(n100), .B1(
        \REGISTERS[19][28] ), .B2(n99), .ZN(n1280) );
  AOI22_X1 U1314 ( .A1(\REGISTERS[20][28] ), .A2(n102), .B1(
        \REGISTERS[21][28] ), .B2(n101), .ZN(n1279) );
  AOI22_X1 U1315 ( .A1(\REGISTERS[4][28] ), .A2(n104), .B1(\REGISTERS[2][28] ), 
        .B2(n103), .ZN(n1278) );
  AOI22_X1 U1316 ( .A1(\REGISTERS[26][28] ), .A2(n106), .B1(
        \REGISTERS[27][28] ), .B2(n105), .ZN(n1264) );
  AOI22_X1 U1317 ( .A1(\REGISTERS[28][28] ), .A2(n108), .B1(
        \REGISTERS[29][28] ), .B2(n107), .ZN(n1263) );
  AOI22_X1 U1318 ( .A1(\REGISTERS[30][28] ), .A2(n1492), .B1(
        \REGISTERS[7][28] ), .B2(n109), .ZN(n1262) );
  AOI22_X1 U1319 ( .A1(\REGISTERS[5][28] ), .A2(n1494), .B1(\REGISTERS[3][28] ), .B2(n111), .ZN(n1261) );
  NAND4_X1 U1320 ( .A1(n1264), .A2(n1263), .A3(n1262), .A4(n1261), .ZN(n1276)
         );
  AOI22_X1 U1321 ( .A1(\REGISTERS[9][28] ), .A2(n114), .B1(\REGISTERS[10][28] ), .B2(n113), .ZN(n1268) );
  AOI22_X1 U1322 ( .A1(\REGISTERS[11][28] ), .A2(n116), .B1(
        \REGISTERS[12][28] ), .B2(n115), .ZN(n1267) );
  AOI22_X1 U1323 ( .A1(\REGISTERS[13][28] ), .A2(n118), .B1(
        \REGISTERS[14][28] ), .B2(n117), .ZN(n1266) );
  AOI22_X1 U1324 ( .A1(\REGISTERS[15][28] ), .A2(n120), .B1(
        \REGISTERS[17][28] ), .B2(n119), .ZN(n1265) );
  NAND4_X1 U1325 ( .A1(n1268), .A2(n1267), .A3(n1266), .A4(n1265), .ZN(n1275)
         );
  AOI22_X1 U1326 ( .A1(\REGISTERS[31][28] ), .A2(n1512), .B1(
        \REGISTERS[22][28] ), .B2(n121), .ZN(n1269) );
  OAI21_X1 U1327 ( .B1(n58), .B2(n1514), .A(n1269), .ZN(n1274) );
  AOI22_X1 U1328 ( .A1(\REGISTERS[24][28] ), .A2(n124), .B1(
        \REGISTERS[25][28] ), .B2(n123), .ZN(n1272) );
  AOI22_X1 U1329 ( .A1(\REGISTERS[8][28] ), .A2(n36), .B1(\REGISTERS[23][28] ), 
        .B2(n125), .ZN(n1271) );
  AOI22_X1 U1330 ( .A1(\REGISTERS[16][28] ), .A2(n1520), .B1(
        \REGISTERS[1][28] ), .B2(n37), .ZN(n1270) );
  NAND3_X1 U1331 ( .A1(n1272), .A2(n1271), .A3(n1270), .ZN(n1273) );
  NOR4_X1 U1332 ( .A1(n1276), .A2(n1275), .A3(n1274), .A4(n1273), .ZN(n1277)
         );
  NAND4_X1 U1333 ( .A1(n1280), .A2(n1279), .A3(n1278), .A4(n1277), .ZN(
        OUT2[28]) );
  AOI22_X1 U1334 ( .A1(\REGISTERS[18][29] ), .A2(n100), .B1(
        \REGISTERS[19][29] ), .B2(n99), .ZN(n1300) );
  AOI22_X1 U1335 ( .A1(\REGISTERS[20][29] ), .A2(n102), .B1(
        \REGISTERS[21][29] ), .B2(n101), .ZN(n1299) );
  AOI22_X1 U1336 ( .A1(\REGISTERS[4][29] ), .A2(n104), .B1(\REGISTERS[2][29] ), 
        .B2(n103), .ZN(n1298) );
  AOI22_X1 U1337 ( .A1(\REGISTERS[26][29] ), .A2(n1488), .B1(
        \REGISTERS[27][29] ), .B2(n105), .ZN(n1284) );
  AOI22_X1 U1338 ( .A1(\REGISTERS[28][29] ), .A2(n1490), .B1(
        \REGISTERS[29][29] ), .B2(n107), .ZN(n1283) );
  AOI22_X1 U1339 ( .A1(\REGISTERS[30][29] ), .A2(n1492), .B1(
        \REGISTERS[7][29] ), .B2(n109), .ZN(n1282) );
  AOI22_X1 U1340 ( .A1(\REGISTERS[5][29] ), .A2(n1494), .B1(\REGISTERS[3][29] ), .B2(n111), .ZN(n1281) );
  NAND4_X1 U1341 ( .A1(n1284), .A2(n1283), .A3(n1282), .A4(n1281), .ZN(n1296)
         );
  AOI22_X1 U1342 ( .A1(\REGISTERS[9][29] ), .A2(n1500), .B1(
        \REGISTERS[10][29] ), .B2(n113), .ZN(n1288) );
  AOI22_X1 U1343 ( .A1(\REGISTERS[11][29] ), .A2(n1502), .B1(
        \REGISTERS[12][29] ), .B2(n115), .ZN(n1287) );
  AOI22_X1 U1344 ( .A1(\REGISTERS[13][29] ), .A2(n1504), .B1(
        \REGISTERS[14][29] ), .B2(n117), .ZN(n1286) );
  AOI22_X1 U1345 ( .A1(\REGISTERS[15][29] ), .A2(n1506), .B1(
        \REGISTERS[17][29] ), .B2(n119), .ZN(n1285) );
  NAND4_X1 U1346 ( .A1(n1288), .A2(n1287), .A3(n1286), .A4(n1285), .ZN(n1295)
         );
  AOI22_X1 U1347 ( .A1(\REGISTERS[31][29] ), .A2(n1512), .B1(
        \REGISTERS[22][29] ), .B2(n121), .ZN(n1289) );
  OAI21_X1 U1348 ( .B1(n59), .B2(n1514), .A(n1289), .ZN(n1294) );
  AOI22_X1 U1349 ( .A1(\REGISTERS[24][29] ), .A2(n1516), .B1(
        \REGISTERS[25][29] ), .B2(n123), .ZN(n1292) );
  AOI22_X1 U1350 ( .A1(\REGISTERS[8][29] ), .A2(n36), .B1(\REGISTERS[23][29] ), 
        .B2(n125), .ZN(n1291) );
  AOI22_X1 U1351 ( .A1(\REGISTERS[16][29] ), .A2(n1520), .B1(
        \REGISTERS[1][29] ), .B2(n37), .ZN(n1290) );
  NAND3_X1 U1352 ( .A1(n1292), .A2(n1291), .A3(n1290), .ZN(n1293) );
  NOR4_X1 U1353 ( .A1(n1296), .A2(n1295), .A3(n1294), .A4(n1293), .ZN(n1297)
         );
  NAND4_X1 U1354 ( .A1(n1300), .A2(n1299), .A3(n1298), .A4(n1297), .ZN(
        OUT2[29]) );
  AOI22_X1 U1355 ( .A1(\REGISTERS[18][2] ), .A2(n1482), .B1(\REGISTERS[19][2] ), .B2(n1481), .ZN(n1320) );
  AOI22_X1 U1356 ( .A1(\REGISTERS[20][2] ), .A2(n1484), .B1(\REGISTERS[21][2] ), .B2(n1483), .ZN(n1319) );
  AOI22_X1 U1357 ( .A1(\REGISTERS[4][2] ), .A2(n1486), .B1(\REGISTERS[2][2] ), 
        .B2(n1485), .ZN(n1318) );
  AOI22_X1 U1358 ( .A1(\REGISTERS[26][2] ), .A2(n1488), .B1(\REGISTERS[27][2] ), .B2(n1487), .ZN(n1304) );
  AOI22_X1 U1359 ( .A1(\REGISTERS[28][2] ), .A2(n1490), .B1(\REGISTERS[29][2] ), .B2(n1489), .ZN(n1303) );
  AOI22_X1 U1360 ( .A1(\REGISTERS[30][2] ), .A2(n1492), .B1(\REGISTERS[7][2] ), 
        .B2(n1491), .ZN(n1302) );
  AOI22_X1 U1361 ( .A1(\REGISTERS[5][2] ), .A2(n1494), .B1(\REGISTERS[3][2] ), 
        .B2(n1493), .ZN(n1301) );
  NAND4_X1 U1362 ( .A1(n1304), .A2(n1303), .A3(n1302), .A4(n1301), .ZN(n1316)
         );
  AOI22_X1 U1363 ( .A1(\REGISTERS[9][2] ), .A2(n1500), .B1(\REGISTERS[10][2] ), 
        .B2(n1499), .ZN(n1308) );
  AOI22_X1 U1364 ( .A1(\REGISTERS[11][2] ), .A2(n1502), .B1(\REGISTERS[12][2] ), .B2(n1501), .ZN(n1307) );
  AOI22_X1 U1365 ( .A1(\REGISTERS[13][2] ), .A2(n1504), .B1(\REGISTERS[14][2] ), .B2(n1503), .ZN(n1306) );
  AOI22_X1 U1366 ( .A1(\REGISTERS[15][2] ), .A2(n1506), .B1(\REGISTERS[17][2] ), .B2(n1505), .ZN(n1305) );
  NAND4_X1 U1367 ( .A1(n1308), .A2(n1307), .A3(n1306), .A4(n1305), .ZN(n1315)
         );
  AOI22_X1 U1368 ( .A1(\REGISTERS[31][2] ), .A2(n1512), .B1(\REGISTERS[22][2] ), .B2(n1511), .ZN(n1309) );
  OAI21_X1 U1369 ( .B1(n60), .B2(n1514), .A(n1309), .ZN(n1314) );
  AOI22_X1 U1370 ( .A1(\REGISTERS[24][2] ), .A2(n1516), .B1(\REGISTERS[25][2] ), .B2(n1515), .ZN(n1312) );
  AOI22_X1 U1371 ( .A1(\REGISTERS[8][2] ), .A2(n36), .B1(\REGISTERS[23][2] ), 
        .B2(n1517), .ZN(n1311) );
  AOI22_X1 U1372 ( .A1(\REGISTERS[16][2] ), .A2(n1520), .B1(\REGISTERS[1][2] ), 
        .B2(n37), .ZN(n1310) );
  NAND3_X1 U1373 ( .A1(n1312), .A2(n1311), .A3(n1310), .ZN(n1313) );
  NOR4_X1 U1374 ( .A1(n1316), .A2(n1315), .A3(n1314), .A4(n1313), .ZN(n1317)
         );
  NAND4_X1 U1375 ( .A1(n1320), .A2(n1319), .A3(n1318), .A4(n1317), .ZN(OUT2[2]) );
  AOI22_X1 U1376 ( .A1(\REGISTERS[18][30] ), .A2(n1482), .B1(
        \REGISTERS[19][30] ), .B2(n1481), .ZN(n1340) );
  AOI22_X1 U1377 ( .A1(\REGISTERS[20][30] ), .A2(n1484), .B1(
        \REGISTERS[21][30] ), .B2(n1483), .ZN(n1339) );
  AOI22_X1 U1378 ( .A1(\REGISTERS[4][30] ), .A2(n1486), .B1(\REGISTERS[2][30] ), .B2(n1485), .ZN(n1338) );
  AOI22_X1 U1379 ( .A1(\REGISTERS[26][30] ), .A2(n1488), .B1(
        \REGISTERS[27][30] ), .B2(n1487), .ZN(n1324) );
  AOI22_X1 U1380 ( .A1(\REGISTERS[28][30] ), .A2(n1490), .B1(
        \REGISTERS[29][30] ), .B2(n1489), .ZN(n1323) );
  AOI22_X1 U1381 ( .A1(\REGISTERS[30][30] ), .A2(n1492), .B1(
        \REGISTERS[7][30] ), .B2(n1491), .ZN(n1322) );
  AOI22_X1 U1382 ( .A1(\REGISTERS[5][30] ), .A2(n1494), .B1(\REGISTERS[3][30] ), .B2(n1493), .ZN(n1321) );
  NAND4_X1 U1383 ( .A1(n1324), .A2(n1323), .A3(n1322), .A4(n1321), .ZN(n1336)
         );
  AOI22_X1 U1384 ( .A1(\REGISTERS[9][30] ), .A2(n1500), .B1(
        \REGISTERS[10][30] ), .B2(n1499), .ZN(n1328) );
  AOI22_X1 U1385 ( .A1(\REGISTERS[11][30] ), .A2(n1502), .B1(
        \REGISTERS[12][30] ), .B2(n1501), .ZN(n1327) );
  AOI22_X1 U1386 ( .A1(\REGISTERS[13][30] ), .A2(n1504), .B1(
        \REGISTERS[14][30] ), .B2(n1503), .ZN(n1326) );
  AOI22_X1 U1387 ( .A1(\REGISTERS[15][30] ), .A2(n1506), .B1(
        \REGISTERS[17][30] ), .B2(n1505), .ZN(n1325) );
  NAND4_X1 U1388 ( .A1(n1328), .A2(n1327), .A3(n1326), .A4(n1325), .ZN(n1335)
         );
  AOI22_X1 U1389 ( .A1(\REGISTERS[31][30] ), .A2(n1512), .B1(
        \REGISTERS[22][30] ), .B2(n1511), .ZN(n1329) );
  OAI21_X1 U1390 ( .B1(n61), .B2(n1514), .A(n1329), .ZN(n1334) );
  AOI22_X1 U1391 ( .A1(\REGISTERS[24][30] ), .A2(n1516), .B1(
        \REGISTERS[25][30] ), .B2(n1515), .ZN(n1332) );
  AOI22_X1 U1392 ( .A1(\REGISTERS[8][30] ), .A2(n36), .B1(\REGISTERS[23][30] ), 
        .B2(n1517), .ZN(n1331) );
  AOI22_X1 U1393 ( .A1(\REGISTERS[16][30] ), .A2(n1520), .B1(
        \REGISTERS[1][30] ), .B2(n37), .ZN(n1330) );
  NAND3_X1 U1394 ( .A1(n1332), .A2(n1331), .A3(n1330), .ZN(n1333) );
  NOR4_X1 U1395 ( .A1(n1336), .A2(n1335), .A3(n1334), .A4(n1333), .ZN(n1337)
         );
  NAND4_X1 U1396 ( .A1(n1340), .A2(n1339), .A3(n1338), .A4(n1337), .ZN(
        OUT2[30]) );
  AOI22_X1 U1397 ( .A1(\REGISTERS[18][31] ), .A2(n1482), .B1(
        \REGISTERS[19][31] ), .B2(n1481), .ZN(n1360) );
  AOI22_X1 U1398 ( .A1(\REGISTERS[20][31] ), .A2(n1484), .B1(
        \REGISTERS[21][31] ), .B2(n1483), .ZN(n1359) );
  AOI22_X1 U1399 ( .A1(\REGISTERS[4][31] ), .A2(n1486), .B1(\REGISTERS[2][31] ), .B2(n1485), .ZN(n1358) );
  AOI22_X1 U1400 ( .A1(\REGISTERS[26][31] ), .A2(n1488), .B1(
        \REGISTERS[27][31] ), .B2(n1487), .ZN(n1344) );
  AOI22_X1 U1401 ( .A1(\REGISTERS[28][31] ), .A2(n1490), .B1(
        \REGISTERS[29][31] ), .B2(n1489), .ZN(n1343) );
  AOI22_X1 U1402 ( .A1(\REGISTERS[30][31] ), .A2(n1492), .B1(
        \REGISTERS[7][31] ), .B2(n1491), .ZN(n1342) );
  AOI22_X1 U1403 ( .A1(\REGISTERS[5][31] ), .A2(n1494), .B1(\REGISTERS[3][31] ), .B2(n1493), .ZN(n1341) );
  NAND4_X1 U1404 ( .A1(n1344), .A2(n1343), .A3(n1342), .A4(n1341), .ZN(n1356)
         );
  AOI22_X1 U1405 ( .A1(\REGISTERS[9][31] ), .A2(n1500), .B1(
        \REGISTERS[10][31] ), .B2(n1499), .ZN(n1348) );
  AOI22_X1 U1406 ( .A1(\REGISTERS[11][31] ), .A2(n1502), .B1(
        \REGISTERS[12][31] ), .B2(n1501), .ZN(n1347) );
  AOI22_X1 U1407 ( .A1(\REGISTERS[13][31] ), .A2(n1504), .B1(
        \REGISTERS[14][31] ), .B2(n1503), .ZN(n1346) );
  AOI22_X1 U1408 ( .A1(\REGISTERS[15][31] ), .A2(n1506), .B1(
        \REGISTERS[17][31] ), .B2(n1505), .ZN(n1345) );
  NAND4_X1 U1409 ( .A1(n1348), .A2(n1347), .A3(n1346), .A4(n1345), .ZN(n1355)
         );
  AOI22_X1 U1410 ( .A1(\REGISTERS[31][31] ), .A2(n1512), .B1(
        \REGISTERS[22][31] ), .B2(n1511), .ZN(n1349) );
  OAI21_X1 U1411 ( .B1(n62), .B2(n1514), .A(n1349), .ZN(n1354) );
  AOI22_X1 U1412 ( .A1(\REGISTERS[24][31] ), .A2(n1516), .B1(
        \REGISTERS[25][31] ), .B2(n1515), .ZN(n1352) );
  AOI22_X1 U1413 ( .A1(\REGISTERS[8][31] ), .A2(n36), .B1(\REGISTERS[23][31] ), 
        .B2(n1517), .ZN(n1351) );
  AOI22_X1 U1414 ( .A1(\REGISTERS[16][31] ), .A2(n1520), .B1(
        \REGISTERS[1][31] ), .B2(n37), .ZN(n1350) );
  NAND3_X1 U1415 ( .A1(n1352), .A2(n1351), .A3(n1350), .ZN(n1353) );
  NOR4_X1 U1416 ( .A1(n1356), .A2(n1355), .A3(n1354), .A4(n1353), .ZN(n1357)
         );
  NAND4_X1 U1417 ( .A1(n1360), .A2(n1359), .A3(n1358), .A4(n1357), .ZN(
        OUT2[31]) );
  AOI22_X1 U1418 ( .A1(\REGISTERS[18][3] ), .A2(n1482), .B1(\REGISTERS[19][3] ), .B2(n1481), .ZN(n1380) );
  AOI22_X1 U1419 ( .A1(\REGISTERS[20][3] ), .A2(n1484), .B1(\REGISTERS[21][3] ), .B2(n1483), .ZN(n1379) );
  AOI22_X1 U1420 ( .A1(\REGISTERS[4][3] ), .A2(n1486), .B1(\REGISTERS[2][3] ), 
        .B2(n1485), .ZN(n1378) );
  AOI22_X1 U1421 ( .A1(\REGISTERS[26][3] ), .A2(n1488), .B1(\REGISTERS[27][3] ), .B2(n1487), .ZN(n1364) );
  AOI22_X1 U1422 ( .A1(\REGISTERS[28][3] ), .A2(n1490), .B1(\REGISTERS[29][3] ), .B2(n1489), .ZN(n1363) );
  AOI22_X1 U1423 ( .A1(\REGISTERS[30][3] ), .A2(n1492), .B1(\REGISTERS[7][3] ), 
        .B2(n1491), .ZN(n1362) );
  AOI22_X1 U1424 ( .A1(\REGISTERS[5][3] ), .A2(n1494), .B1(\REGISTERS[3][3] ), 
        .B2(n1493), .ZN(n1361) );
  NAND4_X1 U1425 ( .A1(n1364), .A2(n1363), .A3(n1362), .A4(n1361), .ZN(n1376)
         );
  AOI22_X1 U1426 ( .A1(\REGISTERS[9][3] ), .A2(n1500), .B1(\REGISTERS[10][3] ), 
        .B2(n1499), .ZN(n1368) );
  AOI22_X1 U1427 ( .A1(\REGISTERS[11][3] ), .A2(n1502), .B1(\REGISTERS[12][3] ), .B2(n1501), .ZN(n1367) );
  AOI22_X1 U1428 ( .A1(\REGISTERS[13][3] ), .A2(n1504), .B1(\REGISTERS[14][3] ), .B2(n1503), .ZN(n1366) );
  AOI22_X1 U1429 ( .A1(\REGISTERS[15][3] ), .A2(n1506), .B1(\REGISTERS[17][3] ), .B2(n1505), .ZN(n1365) );
  NAND4_X1 U1430 ( .A1(n1368), .A2(n1367), .A3(n1366), .A4(n1365), .ZN(n1375)
         );
  AOI22_X1 U1431 ( .A1(\REGISTERS[31][3] ), .A2(n1512), .B1(\REGISTERS[22][3] ), .B2(n1511), .ZN(n1369) );
  OAI21_X1 U1432 ( .B1(n63), .B2(n1514), .A(n1369), .ZN(n1374) );
  AOI22_X1 U1433 ( .A1(\REGISTERS[24][3] ), .A2(n1516), .B1(\REGISTERS[25][3] ), .B2(n1515), .ZN(n1372) );
  AOI22_X1 U1434 ( .A1(\REGISTERS[8][3] ), .A2(n1518), .B1(\REGISTERS[23][3] ), 
        .B2(n1517), .ZN(n1371) );
  AOI22_X1 U1435 ( .A1(\REGISTERS[16][3] ), .A2(n1520), .B1(\REGISTERS[1][3] ), 
        .B2(n1519), .ZN(n1370) );
  NAND3_X1 U1436 ( .A1(n1372), .A2(n1371), .A3(n1370), .ZN(n1373) );
  NOR4_X1 U1437 ( .A1(n1376), .A2(n1375), .A3(n1374), .A4(n1373), .ZN(n1377)
         );
  NAND4_X1 U1438 ( .A1(n1380), .A2(n1379), .A3(n1378), .A4(n1377), .ZN(OUT2[3]) );
  AOI22_X1 U1439 ( .A1(\REGISTERS[18][4] ), .A2(n1482), .B1(\REGISTERS[19][4] ), .B2(n1481), .ZN(n1400) );
  AOI22_X1 U1440 ( .A1(\REGISTERS[20][4] ), .A2(n1484), .B1(\REGISTERS[21][4] ), .B2(n1483), .ZN(n1399) );
  AOI22_X1 U1441 ( .A1(\REGISTERS[4][4] ), .A2(n1486), .B1(\REGISTERS[2][4] ), 
        .B2(n1485), .ZN(n1398) );
  AOI22_X1 U1442 ( .A1(\REGISTERS[26][4] ), .A2(n1488), .B1(\REGISTERS[27][4] ), .B2(n1487), .ZN(n1384) );
  AOI22_X1 U1443 ( .A1(\REGISTERS[28][4] ), .A2(n1490), .B1(\REGISTERS[29][4] ), .B2(n1489), .ZN(n1383) );
  AOI22_X1 U1444 ( .A1(\REGISTERS[30][4] ), .A2(n1492), .B1(\REGISTERS[7][4] ), 
        .B2(n1491), .ZN(n1382) );
  AOI22_X1 U1445 ( .A1(\REGISTERS[5][4] ), .A2(n1494), .B1(\REGISTERS[3][4] ), 
        .B2(n1493), .ZN(n1381) );
  NAND4_X1 U1446 ( .A1(n1384), .A2(n1383), .A3(n1382), .A4(n1381), .ZN(n1396)
         );
  AOI22_X1 U1447 ( .A1(\REGISTERS[9][4] ), .A2(n1500), .B1(\REGISTERS[10][4] ), 
        .B2(n1499), .ZN(n1388) );
  AOI22_X1 U1448 ( .A1(\REGISTERS[11][4] ), .A2(n1502), .B1(\REGISTERS[12][4] ), .B2(n1501), .ZN(n1387) );
  AOI22_X1 U1449 ( .A1(\REGISTERS[13][4] ), .A2(n1504), .B1(\REGISTERS[14][4] ), .B2(n1503), .ZN(n1386) );
  AOI22_X1 U1450 ( .A1(\REGISTERS[15][4] ), .A2(n1506), .B1(\REGISTERS[17][4] ), .B2(n1505), .ZN(n1385) );
  NAND4_X1 U1451 ( .A1(n1388), .A2(n1387), .A3(n1386), .A4(n1385), .ZN(n1395)
         );
  AOI22_X1 U1452 ( .A1(\REGISTERS[31][4] ), .A2(n1512), .B1(\REGISTERS[22][4] ), .B2(n1511), .ZN(n1389) );
  OAI21_X1 U1453 ( .B1(n64), .B2(n1514), .A(n1389), .ZN(n1394) );
  AOI22_X1 U1454 ( .A1(\REGISTERS[24][4] ), .A2(n1516), .B1(\REGISTERS[25][4] ), .B2(n1515), .ZN(n1392) );
  AOI22_X1 U1455 ( .A1(\REGISTERS[8][4] ), .A2(n1518), .B1(\REGISTERS[23][4] ), 
        .B2(n1517), .ZN(n1391) );
  AOI22_X1 U1456 ( .A1(\REGISTERS[16][4] ), .A2(n1520), .B1(\REGISTERS[1][4] ), 
        .B2(n1519), .ZN(n1390) );
  NAND3_X1 U1457 ( .A1(n1392), .A2(n1391), .A3(n1390), .ZN(n1393) );
  NOR4_X1 U1458 ( .A1(n1396), .A2(n1395), .A3(n1394), .A4(n1393), .ZN(n1397)
         );
  NAND4_X1 U1459 ( .A1(n1400), .A2(n1399), .A3(n1398), .A4(n1397), .ZN(OUT2[4]) );
  AOI22_X1 U1460 ( .A1(\REGISTERS[18][5] ), .A2(n1482), .B1(\REGISTERS[19][5] ), .B2(n1481), .ZN(n1420) );
  AOI22_X1 U1461 ( .A1(\REGISTERS[20][5] ), .A2(n1484), .B1(\REGISTERS[21][5] ), .B2(n1483), .ZN(n1419) );
  AOI22_X1 U1462 ( .A1(\REGISTERS[4][5] ), .A2(n1486), .B1(\REGISTERS[2][5] ), 
        .B2(n1485), .ZN(n1418) );
  AOI22_X1 U1463 ( .A1(\REGISTERS[26][5] ), .A2(n1488), .B1(\REGISTERS[27][5] ), .B2(n1487), .ZN(n1404) );
  AOI22_X1 U1464 ( .A1(\REGISTERS[28][5] ), .A2(n1490), .B1(\REGISTERS[29][5] ), .B2(n1489), .ZN(n1403) );
  AOI22_X1 U1465 ( .A1(\REGISTERS[30][5] ), .A2(n1492), .B1(\REGISTERS[7][5] ), 
        .B2(n1491), .ZN(n1402) );
  AOI22_X1 U1466 ( .A1(\REGISTERS[5][5] ), .A2(n1494), .B1(\REGISTERS[3][5] ), 
        .B2(n1493), .ZN(n1401) );
  NAND4_X1 U1467 ( .A1(n1404), .A2(n1403), .A3(n1402), .A4(n1401), .ZN(n1416)
         );
  AOI22_X1 U1468 ( .A1(\REGISTERS[9][5] ), .A2(n1500), .B1(\REGISTERS[10][5] ), 
        .B2(n1499), .ZN(n1408) );
  AOI22_X1 U1469 ( .A1(\REGISTERS[11][5] ), .A2(n1502), .B1(\REGISTERS[12][5] ), .B2(n1501), .ZN(n1407) );
  AOI22_X1 U1470 ( .A1(\REGISTERS[13][5] ), .A2(n1504), .B1(\REGISTERS[14][5] ), .B2(n1503), .ZN(n1406) );
  AOI22_X1 U1471 ( .A1(\REGISTERS[15][5] ), .A2(n1506), .B1(\REGISTERS[17][5] ), .B2(n1505), .ZN(n1405) );
  NAND4_X1 U1472 ( .A1(n1408), .A2(n1407), .A3(n1406), .A4(n1405), .ZN(n1415)
         );
  AOI22_X1 U1473 ( .A1(\REGISTERS[31][5] ), .A2(n122), .B1(\REGISTERS[22][5] ), 
        .B2(n1511), .ZN(n1409) );
  OAI21_X1 U1474 ( .B1(n65), .B2(n1514), .A(n1409), .ZN(n1414) );
  AOI22_X1 U1475 ( .A1(\REGISTERS[24][5] ), .A2(n1516), .B1(\REGISTERS[25][5] ), .B2(n1515), .ZN(n1412) );
  AOI22_X1 U1476 ( .A1(\REGISTERS[8][5] ), .A2(n1518), .B1(\REGISTERS[23][5] ), 
        .B2(n1517), .ZN(n1411) );
  AOI22_X1 U1477 ( .A1(\REGISTERS[16][5] ), .A2(n1520), .B1(\REGISTERS[1][5] ), 
        .B2(n1519), .ZN(n1410) );
  NAND3_X1 U1478 ( .A1(n1412), .A2(n1411), .A3(n1410), .ZN(n1413) );
  NOR4_X1 U1479 ( .A1(n1416), .A2(n1415), .A3(n1414), .A4(n1413), .ZN(n1417)
         );
  NAND4_X1 U1480 ( .A1(n1420), .A2(n1419), .A3(n1418), .A4(n1417), .ZN(OUT2[5]) );
  AOI22_X1 U1481 ( .A1(\REGISTERS[18][6] ), .A2(n1482), .B1(\REGISTERS[19][6] ), .B2(n1481), .ZN(n1440) );
  AOI22_X1 U1482 ( .A1(\REGISTERS[20][6] ), .A2(n1484), .B1(\REGISTERS[21][6] ), .B2(n1483), .ZN(n1439) );
  AOI22_X1 U1483 ( .A1(\REGISTERS[4][6] ), .A2(n1486), .B1(\REGISTERS[2][6] ), 
        .B2(n1485), .ZN(n1438) );
  AOI22_X1 U1484 ( .A1(\REGISTERS[26][6] ), .A2(n1488), .B1(\REGISTERS[27][6] ), .B2(n1487), .ZN(n1424) );
  AOI22_X1 U1485 ( .A1(\REGISTERS[28][6] ), .A2(n1490), .B1(\REGISTERS[29][6] ), .B2(n1489), .ZN(n1423) );
  AOI22_X1 U1486 ( .A1(\REGISTERS[30][6] ), .A2(n1492), .B1(\REGISTERS[7][6] ), 
        .B2(n1491), .ZN(n1422) );
  AOI22_X1 U1487 ( .A1(\REGISTERS[5][6] ), .A2(n1494), .B1(\REGISTERS[3][6] ), 
        .B2(n1493), .ZN(n1421) );
  NAND4_X1 U1488 ( .A1(n1424), .A2(n1423), .A3(n1422), .A4(n1421), .ZN(n1436)
         );
  AOI22_X1 U1489 ( .A1(\REGISTERS[9][6] ), .A2(n1500), .B1(\REGISTERS[10][6] ), 
        .B2(n1499), .ZN(n1428) );
  AOI22_X1 U1490 ( .A1(\REGISTERS[11][6] ), .A2(n1502), .B1(\REGISTERS[12][6] ), .B2(n1501), .ZN(n1427) );
  AOI22_X1 U1491 ( .A1(\REGISTERS[13][6] ), .A2(n1504), .B1(\REGISTERS[14][6] ), .B2(n1503), .ZN(n1426) );
  AOI22_X1 U1492 ( .A1(\REGISTERS[15][6] ), .A2(n1506), .B1(\REGISTERS[17][6] ), .B2(n1505), .ZN(n1425) );
  NAND4_X1 U1493 ( .A1(n1428), .A2(n1427), .A3(n1426), .A4(n1425), .ZN(n1435)
         );
  AOI22_X1 U1494 ( .A1(\REGISTERS[31][6] ), .A2(n122), .B1(\REGISTERS[22][6] ), 
        .B2(n1511), .ZN(n1429) );
  OAI21_X1 U1495 ( .B1(n66), .B2(n1514), .A(n1429), .ZN(n1434) );
  AOI22_X1 U1496 ( .A1(\REGISTERS[24][6] ), .A2(n1516), .B1(\REGISTERS[25][6] ), .B2(n1515), .ZN(n1432) );
  AOI22_X1 U1497 ( .A1(\REGISTERS[8][6] ), .A2(n1518), .B1(\REGISTERS[23][6] ), 
        .B2(n1517), .ZN(n1431) );
  AOI22_X1 U1498 ( .A1(\REGISTERS[16][6] ), .A2(n1520), .B1(\REGISTERS[1][6] ), 
        .B2(n37), .ZN(n1430) );
  NAND3_X1 U1499 ( .A1(n1432), .A2(n1431), .A3(n1430), .ZN(n1433) );
  NOR4_X1 U1500 ( .A1(n1436), .A2(n1435), .A3(n1434), .A4(n1433), .ZN(n1437)
         );
  NAND4_X1 U1501 ( .A1(n1440), .A2(n1439), .A3(n1438), .A4(n1437), .ZN(OUT2[6]) );
  AOI22_X1 U1502 ( .A1(\REGISTERS[18][7] ), .A2(n1482), .B1(\REGISTERS[19][7] ), .B2(n1481), .ZN(n1460) );
  AOI22_X1 U1503 ( .A1(\REGISTERS[20][7] ), .A2(n1484), .B1(\REGISTERS[21][7] ), .B2(n1483), .ZN(n1459) );
  AOI22_X1 U1504 ( .A1(\REGISTERS[4][7] ), .A2(n1486), .B1(\REGISTERS[2][7] ), 
        .B2(n1485), .ZN(n1458) );
  AOI22_X1 U1505 ( .A1(\REGISTERS[26][7] ), .A2(n1488), .B1(\REGISTERS[27][7] ), .B2(n105), .ZN(n1444) );
  AOI22_X1 U1506 ( .A1(\REGISTERS[28][7] ), .A2(n1490), .B1(\REGISTERS[29][7] ), .B2(n107), .ZN(n1443) );
  AOI22_X1 U1507 ( .A1(\REGISTERS[30][7] ), .A2(n1492), .B1(\REGISTERS[7][7] ), 
        .B2(n109), .ZN(n1442) );
  AOI22_X1 U1508 ( .A1(\REGISTERS[5][7] ), .A2(n112), .B1(\REGISTERS[3][7] ), 
        .B2(n111), .ZN(n1441) );
  NAND4_X1 U1509 ( .A1(n1444), .A2(n1443), .A3(n1442), .A4(n1441), .ZN(n1456)
         );
  AOI22_X1 U1510 ( .A1(\REGISTERS[9][7] ), .A2(n1500), .B1(\REGISTERS[10][7] ), 
        .B2(n1499), .ZN(n1448) );
  AOI22_X1 U1511 ( .A1(\REGISTERS[11][7] ), .A2(n1502), .B1(\REGISTERS[12][7] ), .B2(n1501), .ZN(n1447) );
  AOI22_X1 U1512 ( .A1(\REGISTERS[13][7] ), .A2(n1504), .B1(\REGISTERS[14][7] ), .B2(n1503), .ZN(n1446) );
  AOI22_X1 U1513 ( .A1(\REGISTERS[15][7] ), .A2(n1506), .B1(\REGISTERS[17][7] ), .B2(n1505), .ZN(n1445) );
  NAND4_X1 U1514 ( .A1(n1448), .A2(n1447), .A3(n1446), .A4(n1445), .ZN(n1455)
         );
  AOI22_X1 U1515 ( .A1(\REGISTERS[31][7] ), .A2(n1512), .B1(\REGISTERS[22][7] ), .B2(n1511), .ZN(n1449) );
  OAI21_X1 U1516 ( .B1(n67), .B2(n1514), .A(n1449), .ZN(n1454) );
  AOI22_X1 U1517 ( .A1(\REGISTERS[24][7] ), .A2(n1516), .B1(\REGISTERS[25][7] ), .B2(n123), .ZN(n1452) );
  AOI22_X1 U1518 ( .A1(\REGISTERS[8][7] ), .A2(n1518), .B1(\REGISTERS[23][7] ), 
        .B2(n1517), .ZN(n1451) );
  AOI22_X1 U1519 ( .A1(\REGISTERS[16][7] ), .A2(n1520), .B1(\REGISTERS[1][7] ), 
        .B2(n37), .ZN(n1450) );
  NAND3_X1 U1520 ( .A1(n1452), .A2(n1451), .A3(n1450), .ZN(n1453) );
  NOR4_X1 U1521 ( .A1(n1456), .A2(n1455), .A3(n1454), .A4(n1453), .ZN(n1457)
         );
  NAND4_X1 U1522 ( .A1(n1460), .A2(n1459), .A3(n1458), .A4(n1457), .ZN(OUT2[7]) );
  AOI22_X1 U1523 ( .A1(\REGISTERS[18][8] ), .A2(n100), .B1(\REGISTERS[19][8] ), 
        .B2(n99), .ZN(n1480) );
  AOI22_X1 U1524 ( .A1(\REGISTERS[20][8] ), .A2(n102), .B1(\REGISTERS[21][8] ), 
        .B2(n101), .ZN(n1479) );
  AOI22_X1 U1525 ( .A1(\REGISTERS[4][8] ), .A2(n104), .B1(\REGISTERS[2][8] ), 
        .B2(n103), .ZN(n1478) );
  AOI22_X1 U1526 ( .A1(\REGISTERS[26][8] ), .A2(n1488), .B1(\REGISTERS[27][8] ), .B2(n105), .ZN(n1464) );
  AOI22_X1 U1527 ( .A1(\REGISTERS[28][8] ), .A2(n1490), .B1(\REGISTERS[29][8] ), .B2(n107), .ZN(n1463) );
  AOI22_X1 U1528 ( .A1(\REGISTERS[30][8] ), .A2(n110), .B1(\REGISTERS[7][8] ), 
        .B2(n109), .ZN(n1462) );
  AOI22_X1 U1529 ( .A1(\REGISTERS[5][8] ), .A2(n112), .B1(\REGISTERS[3][8] ), 
        .B2(n111), .ZN(n1461) );
  NAND4_X1 U1530 ( .A1(n1464), .A2(n1463), .A3(n1462), .A4(n1461), .ZN(n1476)
         );
  AOI22_X1 U1531 ( .A1(\REGISTERS[9][8] ), .A2(n1500), .B1(\REGISTERS[10][8] ), 
        .B2(n1499), .ZN(n1468) );
  AOI22_X1 U1532 ( .A1(\REGISTERS[11][8] ), .A2(n1502), .B1(\REGISTERS[12][8] ), .B2(n1501), .ZN(n1467) );
  AOI22_X1 U1533 ( .A1(\REGISTERS[13][8] ), .A2(n1504), .B1(\REGISTERS[14][8] ), .B2(n1503), .ZN(n1466) );
  AOI22_X1 U1534 ( .A1(\REGISTERS[15][8] ), .A2(n1506), .B1(\REGISTERS[17][8] ), .B2(n1505), .ZN(n1465) );
  NAND4_X1 U1535 ( .A1(n1468), .A2(n1467), .A3(n1466), .A4(n1465), .ZN(n1475)
         );
  AOI22_X1 U1536 ( .A1(\REGISTERS[31][8] ), .A2(n1512), .B1(\REGISTERS[22][8] ), .B2(n1511), .ZN(n1469) );
  OAI21_X1 U1537 ( .B1(n68), .B2(n1514), .A(n1469), .ZN(n1474) );
  AOI22_X1 U1538 ( .A1(\REGISTERS[24][8] ), .A2(n1516), .B1(\REGISTERS[25][8] ), .B2(n123), .ZN(n1472) );
  AOI22_X1 U1539 ( .A1(\REGISTERS[8][8] ), .A2(n36), .B1(\REGISTERS[23][8] ), 
        .B2(n1517), .ZN(n1471) );
  AOI22_X1 U1540 ( .A1(\REGISTERS[16][8] ), .A2(n1520), .B1(\REGISTERS[1][8] ), 
        .B2(n37), .ZN(n1470) );
  NAND3_X1 U1541 ( .A1(n1472), .A2(n1471), .A3(n1470), .ZN(n1473) );
  NOR4_X1 U1542 ( .A1(n1476), .A2(n1475), .A3(n1474), .A4(n1473), .ZN(n1477)
         );
  NAND4_X1 U1543 ( .A1(n1480), .A2(n1479), .A3(n1478), .A4(n1477), .ZN(OUT2[8]) );
  AOI22_X1 U1544 ( .A1(\REGISTERS[18][9] ), .A2(n100), .B1(\REGISTERS[19][9] ), 
        .B2(n99), .ZN(n1531) );
  AOI22_X1 U1545 ( .A1(\REGISTERS[20][9] ), .A2(n102), .B1(\REGISTERS[21][9] ), 
        .B2(n101), .ZN(n1530) );
  AOI22_X1 U1546 ( .A1(\REGISTERS[4][9] ), .A2(n104), .B1(\REGISTERS[2][9] ), 
        .B2(n103), .ZN(n1529) );
  AOI22_X1 U1547 ( .A1(\REGISTERS[26][9] ), .A2(n106), .B1(\REGISTERS[27][9] ), 
        .B2(n105), .ZN(n1498) );
  AOI22_X1 U1548 ( .A1(\REGISTERS[28][9] ), .A2(n108), .B1(\REGISTERS[29][9] ), 
        .B2(n107), .ZN(n1497) );
  AOI22_X1 U1549 ( .A1(\REGISTERS[30][9] ), .A2(n110), .B1(\REGISTERS[7][9] ), 
        .B2(n109), .ZN(n1496) );
  AOI22_X1 U1550 ( .A1(\REGISTERS[5][9] ), .A2(n112), .B1(\REGISTERS[3][9] ), 
        .B2(n111), .ZN(n1495) );
  NAND4_X1 U1551 ( .A1(n1498), .A2(n1497), .A3(n1496), .A4(n1495), .ZN(n1527)
         );
  AOI22_X1 U1552 ( .A1(\REGISTERS[9][9] ), .A2(n114), .B1(\REGISTERS[10][9] ), 
        .B2(n113), .ZN(n1510) );
  AOI22_X1 U1553 ( .A1(\REGISTERS[11][9] ), .A2(n116), .B1(\REGISTERS[12][9] ), 
        .B2(n115), .ZN(n1509) );
  AOI22_X1 U1554 ( .A1(\REGISTERS[13][9] ), .A2(n118), .B1(\REGISTERS[14][9] ), 
        .B2(n117), .ZN(n1508) );
  AOI22_X1 U1555 ( .A1(\REGISTERS[15][9] ), .A2(n120), .B1(\REGISTERS[17][9] ), 
        .B2(n119), .ZN(n1507) );
  NAND4_X1 U1556 ( .A1(n1510), .A2(n1509), .A3(n1508), .A4(n1507), .ZN(n1526)
         );
  AOI22_X1 U1557 ( .A1(\REGISTERS[31][9] ), .A2(n1512), .B1(\REGISTERS[22][9] ), .B2(n121), .ZN(n1513) );
  OAI21_X1 U1558 ( .B1(n69), .B2(n1514), .A(n1513), .ZN(n1525) );
  AOI22_X1 U1559 ( .A1(\REGISTERS[24][9] ), .A2(n124), .B1(\REGISTERS[25][9] ), 
        .B2(n123), .ZN(n1523) );
  AOI22_X1 U1560 ( .A1(\REGISTERS[8][9] ), .A2(n36), .B1(\REGISTERS[23][9] ), 
        .B2(n125), .ZN(n1522) );
  AOI22_X1 U1561 ( .A1(\REGISTERS[16][9] ), .A2(n1520), .B1(\REGISTERS[1][9] ), 
        .B2(n37), .ZN(n1521) );
  NAND3_X1 U1562 ( .A1(n1523), .A2(n1522), .A3(n1521), .ZN(n1524) );
  NOR4_X1 U1563 ( .A1(n1527), .A2(n1526), .A3(n1525), .A4(n1524), .ZN(n1528)
         );
  NAND4_X1 U1564 ( .A1(n1531), .A2(n1530), .A3(n1529), .A4(n1528), .ZN(OUT2[9]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_reg_N32_9 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18782, net18784, net18786, net18787, net18790, net18793;
  assign net18782 = EN;
  assign net18784 = CLK;
  assign ENCLK = net18786;
  assign net18793 = TE;

  DLL_X1 latch ( .D(net18787), .GN(net18784), .Q(net18790) );
  AND2_X1 main_gate ( .A1(net18790), .A2(net18784), .ZN(net18786) );
  OR2_X1 test_or ( .A1(net18782), .A2(net18793), .ZN(net18787) );
endmodule


module reg_N32_9 ( D, EN, CLK, RST, \Q[31] , \Q[30] , \Q[29] , \Q[28] , 
        \Q[27] , \Q[26] , \Q[25] , \Q[24] , \Q[23] , \Q[22] , \Q[21] , 
        \Q[20]_BAR , \Q[17] , \Q[15] , \Q[11] , \Q[10] , \Q[9] , \Q[8] , 
        \Q[7] , \Q[6] , \Q[5] , \Q[4] , \Q[3] , \Q[2] , \Q[1] , \Q[0] , 
        \Q[19]_BAR , \Q[18]_BAR , \Q[16]_BAR , \Q[14]_BAR , \Q[13]_BAR , 
        \Q[12]_BAR  );
  input [31:0] D;
  input EN, CLK, RST;
  output \Q[31] , \Q[30] , \Q[29] , \Q[28] , \Q[27] , \Q[26] , \Q[25] ,
         \Q[24] , \Q[23] , \Q[22] , \Q[21] , \Q[20]_BAR , \Q[17] , \Q[15] ,
         \Q[11] , \Q[10] , \Q[9] , \Q[8] , \Q[7] , \Q[6] , \Q[5] , \Q[4] ,
         \Q[3] , \Q[2] , \Q[1] , \Q[0] , \Q[19]_BAR , \Q[18]_BAR , \Q[16]_BAR ,
         \Q[14]_BAR , \Q[13]_BAR , \Q[12]_BAR ;
  wire   net18798, n8, n9, n10, n11, n12;
  wire   [31:0] Q;

  SNPS_CLOCK_GATE_HIGH_reg_N32_9 clk_gate_Q_reg ( .CLK(CLK), .EN(EN), .ENCLK(
        net18798), .TE(1'b0) );
  DFFR_X1 \Q_reg[31]  ( .D(D[31]), .CK(net18798), .RN(RST), .Q(Q[31]) );
  DFFR_X1 \Q_reg[30]  ( .D(D[30]), .CK(net18798), .RN(RST), .Q(Q[30]) );
  DFFR_X1 \Q_reg[29]  ( .D(D[29]), .CK(net18798), .RN(RST), .Q(Q[29]) );
  DFFR_X1 \Q_reg[28]  ( .D(D[28]), .CK(net18798), .RN(RST), .Q(Q[28]) );
  DFFR_X1 \Q_reg[27]  ( .D(D[27]), .CK(net18798), .RN(RST), .Q(Q[27]) );
  DFFR_X1 \Q_reg[26]  ( .D(D[26]), .CK(net18798), .RN(RST), .Q(Q[26]) );
  DFFR_X1 \Q_reg[25]  ( .D(D[25]), .CK(net18798), .RN(RST), .Q(Q[25]) );
  DFFR_X1 \Q_reg[24]  ( .D(D[24]), .CK(net18798), .RN(RST), .Q(Q[24]) );
  DFFR_X1 \Q_reg[23]  ( .D(D[23]), .CK(net18798), .RN(RST), .Q(Q[23]) );
  DFFR_X1 \Q_reg[22]  ( .D(D[22]), .CK(net18798), .RN(RST), .Q(Q[22]) );
  DFFR_X1 \Q_reg[21]  ( .D(D[21]), .CK(net18798), .RN(RST), .Q(Q[21]) );
  DFFR_X1 \Q_reg[20]  ( .D(D[20]), .CK(net18798), .RN(RST), .QN(\Q[20]_BAR )
         );
  DFFR_X1 \Q_reg[19]  ( .D(D[19]), .CK(net18798), .RN(RST), .QN(\Q[19]_BAR )
         );
  DFFR_X1 \Q_reg[18]  ( .D(D[18]), .CK(net18798), .RN(RST), .QN(\Q[18]_BAR )
         );
  DFFR_X1 \Q_reg[17]  ( .D(D[17]), .CK(net18798), .RN(RST), .Q(Q[17]) );
  DFFR_X1 \Q_reg[16]  ( .D(D[16]), .CK(net18798), .RN(RST), .QN(\Q[16]_BAR )
         );
  DFFR_X1 \Q_reg[13]  ( .D(D[13]), .CK(net18798), .RN(RST), .QN(\Q[13]_BAR )
         );
  DFFR_X2 \Q_reg[4]  ( .D(D[4]), .CK(net18798), .RN(RST), .Q(Q[4]) );
  DFFR_X1 \Q_reg[2]  ( .D(D[2]), .CK(net18798), .RN(RST), .Q(Q[2]) );
  DFFR_X2 \Q_reg[6]  ( .D(D[6]), .CK(net18798), .RN(RST), .Q(Q[6]) );
  DFFR_X1 \Q_reg[7]  ( .D(D[7]), .CK(net18798), .RN(RST), .Q(Q[7]) );
  DFFR_X1 \Q_reg[8]  ( .D(D[8]), .CK(net18798), .RN(RST), .Q(Q[8]) );
  DFFR_X1 \Q_reg[10]  ( .D(D[10]), .CK(net18798), .RN(RST), .Q(Q[10]) );
  DFFR_X1 \Q_reg[3]  ( .D(D[3]), .CK(net18798), .RN(RST), .Q(Q[3]) );
  DFFS_X1 \Q_reg[1]  ( .D(n10), .CK(net18798), .SN(RST), .QN(Q[1]) );
  DFFS_X1 \Q_reg[0]  ( .D(n11), .CK(net18798), .SN(RST), .QN(Q[0]) );
  DFFS_X1 \Q_reg[12]  ( .D(n9), .CK(net18798), .SN(RST), .Q(\Q[12]_BAR ) );
  DFFS_X1 \Q_reg[14]  ( .D(n8), .CK(net18798), .SN(RST), .Q(\Q[14]_BAR ) );
  DFFR_X2 \Q_reg[9]  ( .D(D[9]), .CK(net18798), .RN(RST), .Q(Q[9]) );
  DFFS_X2 \Q_reg[5]  ( .D(n12), .CK(net18798), .SN(RST), .QN(Q[5]) );
  DFFR_X2 \Q_reg[15]  ( .D(D[15]), .CK(net18798), .RN(RST), .Q(Q[15]) );
  DFFR_X1 \Q_reg[11]  ( .D(D[11]), .CK(net18798), .RN(RST), .Q(Q[11]) );
  INV_X1 U2 ( .A(D[14]), .ZN(n8) );
  INV_X1 U3 ( .A(D[12]), .ZN(n9) );
  INV_X1 U4 ( .A(D[0]), .ZN(n11) );
  INV_X1 U5 ( .A(D[1]), .ZN(n10) );
  INV_X1 U6 ( .A(D[5]), .ZN(n12) );
endmodule


module SNPS_CLOCK_GATE_HIGH_reg_N32_8 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18782, net18784, net18786, net18787, net18790, net18793;
  assign net18782 = EN;
  assign net18784 = CLK;
  assign ENCLK = net18786;
  assign net18793 = TE;

  DLL_X1 latch ( .D(net18787), .GN(net18784), .Q(net18790) );
  AND2_X1 main_gate ( .A1(net18790), .A2(net18784), .ZN(net18786) );
  OR2_X1 test_or ( .A1(net18782), .A2(net18793), .ZN(net18787) );
endmodule


module reg_N32_8 ( D, Q, EN, CLK, RST );
  input [31:0] D;
  output [31:0] Q;
  input EN, CLK, RST;
  wire   net18798;

  SNPS_CLOCK_GATE_HIGH_reg_N32_8 clk_gate_Q_reg ( .CLK(CLK), .EN(EN), .ENCLK(
        net18798), .TE(1'b0) );
  DFFR_X1 \Q_reg[31]  ( .D(D[31]), .CK(net18798), .RN(RST), .Q(Q[31]) );
  DFFR_X1 \Q_reg[30]  ( .D(D[30]), .CK(net18798), .RN(RST), .Q(Q[30]) );
  DFFR_X1 \Q_reg[29]  ( .D(D[29]), .CK(net18798), .RN(RST), .Q(Q[29]) );
  DFFR_X1 \Q_reg[28]  ( .D(D[28]), .CK(net18798), .RN(RST), .Q(Q[28]) );
  DFFR_X1 \Q_reg[27]  ( .D(D[27]), .CK(net18798), .RN(RST), .Q(Q[27]) );
  DFFR_X1 \Q_reg[26]  ( .D(D[26]), .CK(net18798), .RN(RST), .Q(Q[26]) );
  DFFR_X1 \Q_reg[25]  ( .D(D[25]), .CK(net18798), .RN(RST), .Q(Q[25]) );
  DFFR_X1 \Q_reg[24]  ( .D(D[24]), .CK(net18798), .RN(RST), .Q(Q[24]) );
  DFFR_X1 \Q_reg[23]  ( .D(D[23]), .CK(net18798), .RN(RST), .Q(Q[23]) );
  DFFR_X1 \Q_reg[22]  ( .D(D[22]), .CK(net18798), .RN(RST), .Q(Q[22]) );
  DFFR_X1 \Q_reg[21]  ( .D(D[21]), .CK(net18798), .RN(RST), .Q(Q[21]) );
  DFFR_X1 \Q_reg[20]  ( .D(D[20]), .CK(net18798), .RN(RST), .Q(Q[20]) );
  DFFR_X1 \Q_reg[19]  ( .D(D[19]), .CK(net18798), .RN(RST), .Q(Q[19]) );
  DFFR_X1 \Q_reg[18]  ( .D(D[18]), .CK(net18798), .RN(RST), .Q(Q[18]) );
  DFFR_X1 \Q_reg[17]  ( .D(D[17]), .CK(net18798), .RN(RST), .Q(Q[17]) );
  DFFR_X1 \Q_reg[16]  ( .D(D[16]), .CK(net18798), .RN(RST), .Q(Q[16]) );
  DFFR_X1 \Q_reg[15]  ( .D(D[15]), .CK(net18798), .RN(RST), .Q(Q[15]) );
  DFFR_X1 \Q_reg[14]  ( .D(D[14]), .CK(net18798), .RN(RST), .Q(Q[14]) );
  DFFR_X1 \Q_reg[13]  ( .D(D[13]), .CK(net18798), .RN(RST), .Q(Q[13]) );
  DFFR_X1 \Q_reg[12]  ( .D(D[12]), .CK(net18798), .RN(RST), .Q(Q[12]) );
  DFFR_X1 \Q_reg[11]  ( .D(D[11]), .CK(net18798), .RN(RST), .Q(Q[11]) );
  DFFR_X1 \Q_reg[10]  ( .D(D[10]), .CK(net18798), .RN(RST), .Q(Q[10]) );
  DFFR_X1 \Q_reg[9]  ( .D(D[9]), .CK(net18798), .RN(RST), .Q(Q[9]) );
  DFFR_X1 \Q_reg[8]  ( .D(D[8]), .CK(net18798), .RN(RST), .Q(Q[8]) );
  DFFR_X1 \Q_reg[7]  ( .D(D[7]), .CK(net18798), .RN(RST), .Q(Q[7]) );
  DFFR_X1 \Q_reg[6]  ( .D(D[6]), .CK(net18798), .RN(RST), .Q(Q[6]) );
  DFFR_X1 \Q_reg[5]  ( .D(D[5]), .CK(net18798), .RN(RST), .Q(Q[5]) );
  DFFR_X1 \Q_reg[4]  ( .D(D[4]), .CK(net18798), .RN(RST), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(D[3]), .CK(net18798), .RN(RST), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(D[2]), .CK(net18798), .RN(RST), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(D[1]), .CK(net18798), .RN(RST), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(D[0]), .CK(net18798), .RN(RST), .Q(Q[0]) );
endmodule


module MUX_2to1_N32_8 ( IN0, IN1, SEL, Y );
  input [31:0] IN0;
  input [31:0] IN1;
  output [31:0] Y;
  input SEL;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12;
  assign Y[15] = IN0[15];
  assign Y[14] = IN0[14];
  assign Y[13] = IN0[13];
  assign Y[12] = IN0[12];
  assign Y[11] = IN0[11];
  assign Y[10] = IN0[10];
  assign Y[9] = IN0[9];
  assign Y[8] = IN0[8];
  assign Y[7] = IN0[7];
  assign Y[6] = IN0[6];
  assign Y[5] = IN0[5];
  assign Y[4] = IN0[4];
  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];
  assign Y[25] = Y[31];
  assign Y[26] = Y[31];
  assign Y[27] = Y[31];
  assign Y[28] = Y[31];
  assign Y[29] = Y[31];
  assign Y[30] = Y[31];

  NAND2_X2 U1 ( .A1(n12), .A2(n11), .ZN(Y[31]) );
  NAND2_X1 U2 ( .A1(IN0[16]), .A2(n1), .ZN(n12) );
  INV_X1 U3 ( .A(SEL), .ZN(n1) );
  NAND2_X1 U4 ( .A1(SEL), .A2(IN1[16]), .ZN(n2) );
  NAND2_X1 U5 ( .A1(n12), .A2(n2), .ZN(Y[16]) );
  NAND2_X1 U6 ( .A1(SEL), .A2(IN1[17]), .ZN(n3) );
  NAND2_X1 U7 ( .A1(n12), .A2(n3), .ZN(Y[17]) );
  NAND2_X1 U8 ( .A1(SEL), .A2(IN1[18]), .ZN(n4) );
  NAND2_X1 U9 ( .A1(n12), .A2(n4), .ZN(Y[18]) );
  NAND2_X1 U10 ( .A1(SEL), .A2(IN1[19]), .ZN(n5) );
  NAND2_X1 U11 ( .A1(n12), .A2(n5), .ZN(Y[19]) );
  NAND2_X1 U12 ( .A1(SEL), .A2(IN1[20]), .ZN(n6) );
  NAND2_X1 U13 ( .A1(n12), .A2(n6), .ZN(Y[20]) );
  NAND2_X1 U14 ( .A1(SEL), .A2(IN1[21]), .ZN(n7) );
  NAND2_X1 U15 ( .A1(n12), .A2(n7), .ZN(Y[21]) );
  NAND2_X1 U16 ( .A1(SEL), .A2(IN1[22]), .ZN(n8) );
  NAND2_X1 U17 ( .A1(n12), .A2(n8), .ZN(Y[22]) );
  NAND2_X1 U18 ( .A1(SEL), .A2(IN1[23]), .ZN(n9) );
  NAND2_X1 U19 ( .A1(n12), .A2(n9), .ZN(Y[23]) );
  NAND2_X1 U20 ( .A1(SEL), .A2(IN1[24]), .ZN(n10) );
  NAND2_X1 U21 ( .A1(n12), .A2(n10), .ZN(Y[24]) );
  NAND2_X1 U22 ( .A1(SEL), .A2(IN1[25]), .ZN(n11) );
endmodule


module SNPS_CLOCK_GATE_HIGH_reg_N32_7 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18782, net18784, net18786, net18787, net18790, net18793;
  assign net18782 = EN;
  assign net18784 = CLK;
  assign ENCLK = net18786;
  assign net18793 = TE;

  DLL_X1 latch ( .D(net18787), .GN(net18784), .Q(net18790) );
  AND2_X1 main_gate ( .A1(net18790), .A2(net18784), .ZN(net18786) );
  OR2_X1 test_or ( .A1(net18782), .A2(net18793), .ZN(net18787) );
endmodule


module reg_N32_7 ( D, Q, EN, CLK, RST );
  input [31:0] D;
  output [31:0] Q;
  input EN, CLK, RST;
  wire   net18798;

  SNPS_CLOCK_GATE_HIGH_reg_N32_7 clk_gate_Q_reg ( .CLK(CLK), .EN(EN), .ENCLK(
        net18798), .TE(1'b0) );
  DFFR_X1 \Q_reg[31]  ( .D(D[31]), .CK(net18798), .RN(RST), .Q(Q[31]) );
  DFFR_X1 \Q_reg[30]  ( .D(D[30]), .CK(net18798), .RN(RST), .Q(Q[30]) );
  DFFR_X1 \Q_reg[29]  ( .D(D[29]), .CK(net18798), .RN(RST), .Q(Q[29]) );
  DFFR_X1 \Q_reg[28]  ( .D(D[28]), .CK(net18798), .RN(RST), .Q(Q[28]) );
  DFFR_X1 \Q_reg[27]  ( .D(D[27]), .CK(net18798), .RN(RST), .Q(Q[27]) );
  DFFR_X1 \Q_reg[26]  ( .D(D[26]), .CK(net18798), .RN(RST), .Q(Q[26]) );
  DFFR_X1 \Q_reg[25]  ( .D(D[25]), .CK(net18798), .RN(RST), .Q(Q[25]) );
  DFFR_X1 \Q_reg[24]  ( .D(D[24]), .CK(net18798), .RN(RST), .Q(Q[24]) );
  DFFR_X1 \Q_reg[23]  ( .D(D[23]), .CK(net18798), .RN(RST), .Q(Q[23]) );
  DFFR_X1 \Q_reg[22]  ( .D(D[22]), .CK(net18798), .RN(RST), .Q(Q[22]) );
  DFFR_X1 \Q_reg[21]  ( .D(D[21]), .CK(net18798), .RN(RST), .Q(Q[21]) );
  DFFR_X1 \Q_reg[20]  ( .D(D[20]), .CK(net18798), .RN(RST), .Q(Q[20]) );
  DFFR_X1 \Q_reg[19]  ( .D(D[19]), .CK(net18798), .RN(RST), .Q(Q[19]) );
  DFFR_X1 \Q_reg[18]  ( .D(D[18]), .CK(net18798), .RN(RST), .Q(Q[18]) );
  DFFR_X1 \Q_reg[17]  ( .D(D[17]), .CK(net18798), .RN(RST), .Q(Q[17]) );
  DFFR_X1 \Q_reg[16]  ( .D(D[16]), .CK(net18798), .RN(RST), .Q(Q[16]) );
  DFFR_X1 \Q_reg[15]  ( .D(D[15]), .CK(net18798), .RN(RST), .Q(Q[15]) );
  DFFR_X1 \Q_reg[14]  ( .D(D[14]), .CK(net18798), .RN(RST), .Q(Q[14]) );
  DFFR_X1 \Q_reg[13]  ( .D(D[13]), .CK(net18798), .RN(RST), .Q(Q[13]) );
  DFFR_X1 \Q_reg[12]  ( .D(D[12]), .CK(net18798), .RN(RST), .Q(Q[12]) );
  DFFR_X1 \Q_reg[11]  ( .D(D[11]), .CK(net18798), .RN(RST), .Q(Q[11]) );
  DFFR_X1 \Q_reg[10]  ( .D(D[10]), .CK(net18798), .RN(RST), .Q(Q[10]) );
  DFFR_X1 \Q_reg[9]  ( .D(D[9]), .CK(net18798), .RN(RST), .Q(Q[9]) );
  DFFR_X1 \Q_reg[8]  ( .D(D[8]), .CK(net18798), .RN(RST), .Q(Q[8]) );
  DFFR_X1 \Q_reg[7]  ( .D(D[7]), .CK(net18798), .RN(RST), .Q(Q[7]) );
  DFFR_X1 \Q_reg[6]  ( .D(D[6]), .CK(net18798), .RN(RST), .Q(Q[6]) );
  DFFR_X1 \Q_reg[5]  ( .D(D[5]), .CK(net18798), .RN(RST), .Q(Q[5]) );
  DFFR_X1 \Q_reg[4]  ( .D(D[4]), .CK(net18798), .RN(RST), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(D[3]), .CK(net18798), .RN(RST), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(D[2]), .CK(net18798), .RN(RST), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(D[1]), .CK(net18798), .RN(RST), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(D[0]), .CK(net18798), .RN(RST), .Q(Q[0]) );
endmodule


module MUX_2to1_N32_7 ( IN0, IN1, SEL, Y );
  input [31:0] IN0;
  input [31:0] IN1;
  output [31:0] Y;
  input SEL;
  wire   n1, n2;

  BUF_X1 U1 ( .A(SEL), .Z(n1) );
  BUF_X1 U2 ( .A(SEL), .Z(n2) );
  MUX2_X1 U3 ( .A(IN0[0]), .B(IN1[0]), .S(n1), .Z(Y[0]) );
  MUX2_X1 U4 ( .A(IN0[10]), .B(IN1[10]), .S(n1), .Z(Y[10]) );
  MUX2_X1 U5 ( .A(IN0[11]), .B(IN1[11]), .S(n1), .Z(Y[11]) );
  MUX2_X1 U6 ( .A(IN0[12]), .B(IN1[12]), .S(n1), .Z(Y[12]) );
  MUX2_X1 U7 ( .A(IN0[13]), .B(IN1[13]), .S(n1), .Z(Y[13]) );
  MUX2_X1 U8 ( .A(IN0[14]), .B(IN1[14]), .S(n1), .Z(Y[14]) );
  MUX2_X1 U9 ( .A(IN0[15]), .B(IN1[15]), .S(n1), .Z(Y[15]) );
  MUX2_X1 U10 ( .A(IN0[16]), .B(IN1[16]), .S(n1), .Z(Y[16]) );
  MUX2_X1 U11 ( .A(IN0[17]), .B(IN1[17]), .S(n1), .Z(Y[17]) );
  MUX2_X1 U12 ( .A(IN0[18]), .B(IN1[18]), .S(n1), .Z(Y[18]) );
  MUX2_X1 U13 ( .A(IN0[19]), .B(IN1[19]), .S(n1), .Z(Y[19]) );
  MUX2_X1 U14 ( .A(IN0[1]), .B(IN1[1]), .S(n2), .Z(Y[1]) );
  MUX2_X1 U15 ( .A(IN0[20]), .B(IN1[20]), .S(n2), .Z(Y[20]) );
  MUX2_X1 U16 ( .A(IN0[21]), .B(IN1[21]), .S(n2), .Z(Y[21]) );
  MUX2_X1 U17 ( .A(IN0[22]), .B(IN1[22]), .S(n2), .Z(Y[22]) );
  MUX2_X1 U18 ( .A(IN0[23]), .B(IN1[23]), .S(n2), .Z(Y[23]) );
  MUX2_X1 U19 ( .A(IN0[24]), .B(IN1[24]), .S(n2), .Z(Y[24]) );
  MUX2_X1 U20 ( .A(IN0[25]), .B(IN1[25]), .S(n2), .Z(Y[25]) );
  MUX2_X1 U21 ( .A(IN0[26]), .B(IN1[26]), .S(n2), .Z(Y[26]) );
  MUX2_X1 U22 ( .A(IN0[27]), .B(IN1[27]), .S(n2), .Z(Y[27]) );
  MUX2_X1 U23 ( .A(IN0[28]), .B(IN1[28]), .S(n2), .Z(Y[28]) );
  MUX2_X1 U24 ( .A(IN0[29]), .B(IN1[29]), .S(n2), .Z(Y[29]) );
  MUX2_X1 U25 ( .A(IN0[2]), .B(IN1[2]), .S(n2), .Z(Y[2]) );
  MUX2_X1 U26 ( .A(IN0[30]), .B(IN1[30]), .S(n1), .Z(Y[30]) );
  MUX2_X1 U27 ( .A(IN0[31]), .B(IN1[31]), .S(n2), .Z(Y[31]) );
  MUX2_X1 U28 ( .A(IN0[3]), .B(IN1[3]), .S(n1), .Z(Y[3]) );
  MUX2_X1 U29 ( .A(IN0[4]), .B(IN1[4]), .S(SEL), .Z(Y[4]) );
  MUX2_X1 U30 ( .A(IN0[5]), .B(IN1[5]), .S(SEL), .Z(Y[5]) );
  MUX2_X1 U31 ( .A(IN0[6]), .B(IN1[6]), .S(SEL), .Z(Y[6]) );
  MUX2_X1 U32 ( .A(IN0[7]), .B(IN1[7]), .S(SEL), .Z(Y[7]) );
  MUX2_X1 U33 ( .A(IN0[8]), .B(IN1[8]), .S(n2), .Z(Y[8]) );
  MUX2_X1 U34 ( .A(IN0[9]), .B(IN1[9]), .S(n1), .Z(Y[9]) );
endmodule


module MUX_2to1_N32_6 ( IN0, IN1, SEL, Y );
  input [31:0] IN0;
  input [31:0] IN1;
  output [31:0] Y;
  input SEL;
  wire   n1, n2, n3, n4, n5, n6;

  MUX2_X1 U1 ( .A(IN0[5]), .B(IN1[5]), .S(n3), .Z(Y[5]) );
  BUF_X2 U2 ( .A(SEL), .Z(n5) );
  MUX2_X1 U3 ( .A(IN0[3]), .B(IN1[3]), .S(n6), .Z(Y[3]) );
  BUF_X2 U4 ( .A(SEL), .Z(n6) );
  OAI21_X1 U5 ( .B1(n3), .B2(n2), .A(n1), .ZN(Y[2]) );
  NAND2_X1 U6 ( .A1(n6), .A2(IN1[2]), .ZN(n1) );
  INV_X1 U7 ( .A(IN0[2]), .ZN(n2) );
  CLKBUF_X3 U8 ( .A(SEL), .Z(n3) );
  CLKBUF_X3 U9 ( .A(SEL), .Z(n4) );
  MUX2_X1 U10 ( .A(IN0[27]), .B(IN1[27]), .S(n4), .Z(Y[27]) );
  MUX2_X1 U11 ( .A(IN0[9]), .B(IN1[9]), .S(n6), .Z(Y[9]) );
  MUX2_X1 U12 ( .A(IN0[0]), .B(IN1[0]), .S(n6), .Z(Y[0]) );
  MUX2_X1 U13 ( .A(IN0[10]), .B(IN1[10]), .S(n4), .Z(Y[10]) );
  MUX2_X1 U14 ( .A(IN0[11]), .B(IN1[11]), .S(n5), .Z(Y[11]) );
  MUX2_X1 U15 ( .A(IN0[12]), .B(IN1[12]), .S(n3), .Z(Y[12]) );
  MUX2_X1 U16 ( .A(IN0[13]), .B(IN1[13]), .S(n3), .Z(Y[13]) );
  MUX2_X1 U17 ( .A(IN0[14]), .B(IN1[14]), .S(n4), .Z(Y[14]) );
  MUX2_X1 U18 ( .A(IN0[15]), .B(IN1[15]), .S(n3), .Z(Y[15]) );
  MUX2_X1 U19 ( .A(IN0[16]), .B(IN1[16]), .S(n3), .Z(Y[16]) );
  MUX2_X1 U20 ( .A(IN0[17]), .B(IN1[17]), .S(n5), .Z(Y[17]) );
  MUX2_X1 U21 ( .A(IN0[18]), .B(IN1[18]), .S(n3), .Z(Y[18]) );
  MUX2_X1 U22 ( .A(IN0[19]), .B(IN1[19]), .S(n4), .Z(Y[19]) );
  MUX2_X1 U23 ( .A(IN0[1]), .B(IN1[1]), .S(n6), .Z(Y[1]) );
  MUX2_X1 U24 ( .A(IN0[20]), .B(IN1[20]), .S(n5), .Z(Y[20]) );
  MUX2_X1 U25 ( .A(IN0[21]), .B(IN1[21]), .S(n5), .Z(Y[21]) );
  MUX2_X1 U26 ( .A(IN0[22]), .B(IN1[22]), .S(n4), .Z(Y[22]) );
  MUX2_X1 U27 ( .A(IN0[23]), .B(IN1[23]), .S(n3), .Z(Y[23]) );
  MUX2_X1 U28 ( .A(IN0[24]), .B(IN1[24]), .S(n4), .Z(Y[24]) );
  MUX2_X1 U29 ( .A(IN0[25]), .B(IN1[25]), .S(n5), .Z(Y[25]) );
  MUX2_X1 U30 ( .A(IN0[26]), .B(IN1[26]), .S(n4), .Z(Y[26]) );
  MUX2_X1 U31 ( .A(IN0[28]), .B(IN1[28]), .S(n5), .Z(Y[28]) );
  MUX2_X1 U32 ( .A(IN0[29]), .B(IN1[29]), .S(n3), .Z(Y[29]) );
  MUX2_X1 U33 ( .A(IN0[30]), .B(IN1[30]), .S(n4), .Z(Y[30]) );
  MUX2_X1 U34 ( .A(IN0[31]), .B(IN1[31]), .S(n4), .Z(Y[31]) );
  MUX2_X1 U35 ( .A(IN0[4]), .B(IN1[4]), .S(n4), .Z(Y[4]) );
  MUX2_X1 U36 ( .A(IN0[6]), .B(IN1[6]), .S(n5), .Z(Y[6]) );
  MUX2_X1 U37 ( .A(IN0[7]), .B(IN1[7]), .S(n3), .Z(Y[7]) );
  MUX2_X1 U38 ( .A(IN0[8]), .B(IN1[8]), .S(n5), .Z(Y[8]) );
endmodule


module MUX_2to1_N32_4 ( IN0, IN1, SEL, Y );
  input [31:0] IN0;
  input [31:0] IN1;
  output [31:0] Y;
  input SEL;
  wire   n8, n9, n10;

  BUF_X1 U1 ( .A(SEL), .Z(n10) );
  BUF_X1 U2 ( .A(SEL), .Z(n9) );
  BUF_X1 U3 ( .A(SEL), .Z(n8) );
  AND2_X1 U4 ( .A1(n10), .A2(IN1[0]), .ZN(Y[0]) );
  AND2_X1 U5 ( .A1(n10), .A2(IN1[1]), .ZN(Y[1]) );
  AND2_X1 U6 ( .A1(n10), .A2(IN1[2]), .ZN(Y[2]) );
  AND2_X1 U7 ( .A1(n10), .A2(IN1[3]), .ZN(Y[3]) );
  AND2_X1 U8 ( .A1(n10), .A2(IN1[4]), .ZN(Y[4]) );
  AND2_X1 U9 ( .A1(n10), .A2(IN1[5]), .ZN(Y[5]) );
  AND2_X1 U10 ( .A1(n10), .A2(IN1[6]), .ZN(Y[6]) );
  AND2_X1 U11 ( .A1(n10), .A2(IN1[7]), .ZN(Y[7]) );
  AND2_X1 U12 ( .A1(n10), .A2(IN1[8]), .ZN(Y[8]) );
  AND2_X1 U13 ( .A1(n10), .A2(IN1[9]), .ZN(Y[9]) );
  AND2_X1 U14 ( .A1(n10), .A2(IN1[10]), .ZN(Y[10]) );
  AND2_X1 U15 ( .A1(n10), .A2(IN1[11]), .ZN(Y[11]) );
  AND2_X1 U16 ( .A1(n9), .A2(IN1[12]), .ZN(Y[12]) );
  AND2_X1 U17 ( .A1(n9), .A2(IN1[13]), .ZN(Y[13]) );
  AND2_X1 U18 ( .A1(n9), .A2(IN1[14]), .ZN(Y[14]) );
  AND2_X1 U19 ( .A1(n9), .A2(IN1[15]), .ZN(Y[15]) );
  AND2_X1 U20 ( .A1(n9), .A2(IN1[16]), .ZN(Y[16]) );
  AND2_X1 U21 ( .A1(n9), .A2(IN1[17]), .ZN(Y[17]) );
  AND2_X1 U22 ( .A1(n9), .A2(IN1[18]), .ZN(Y[18]) );
  AND2_X1 U23 ( .A1(n9), .A2(IN1[19]), .ZN(Y[19]) );
  AND2_X1 U24 ( .A1(n9), .A2(IN1[20]), .ZN(Y[20]) );
  AND2_X1 U25 ( .A1(n9), .A2(IN1[21]), .ZN(Y[21]) );
  AND2_X1 U26 ( .A1(n8), .A2(IN1[22]), .ZN(Y[22]) );
  AND2_X1 U27 ( .A1(n8), .A2(IN1[23]), .ZN(Y[23]) );
  AND2_X1 U28 ( .A1(n8), .A2(IN1[24]), .ZN(Y[24]) );
  AND2_X1 U29 ( .A1(n8), .A2(IN1[25]), .ZN(Y[25]) );
  AND2_X1 U30 ( .A1(n8), .A2(IN1[26]), .ZN(Y[26]) );
  AND2_X1 U31 ( .A1(n8), .A2(IN1[27]), .ZN(Y[27]) );
  AND2_X1 U32 ( .A1(n8), .A2(IN1[28]), .ZN(Y[28]) );
  AND2_X1 U33 ( .A1(n8), .A2(IN1[29]), .ZN(Y[29]) );
  AND2_X1 U34 ( .A1(n8), .A2(IN1[30]), .ZN(Y[30]) );
  AND2_X1 U35 ( .A1(n8), .A2(IN1[31]), .ZN(Y[31]) );
endmodule


module MUX_2to1_N32_3 ( IN0, IN1, SEL, Y );
  input [31:0] IN0;
  input [31:0] IN1;
  output [31:0] Y;
  input SEL;
  wire   n1, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43;
  assign Y[31] = IN0[31];

  INV_X2 U1 ( .A(n11), .ZN(n1) );
  NAND2_X1 U2 ( .A1(n9), .A2(n12), .ZN(Y[0]) );
  NAND2_X1 U3 ( .A1(n9), .A2(n23), .ZN(Y[1]) );
  CLKBUF_X3 U4 ( .A(n43), .Z(n9) );
  BUF_X1 U5 ( .A(n43), .Z(n10) );
  INV_X1 U6 ( .A(SEL), .ZN(n11) );
  NAND2_X1 U7 ( .A1(IN0[0]), .A2(n11), .ZN(n43) );
  NAND2_X1 U8 ( .A1(n1), .A2(IN1[0]), .ZN(n12) );
  NAND2_X1 U9 ( .A1(n1), .A2(IN1[10]), .ZN(n13) );
  NAND2_X1 U10 ( .A1(n9), .A2(n13), .ZN(Y[10]) );
  NAND2_X1 U11 ( .A1(n1), .A2(IN1[11]), .ZN(n14) );
  NAND2_X1 U12 ( .A1(n9), .A2(n14), .ZN(Y[11]) );
  NAND2_X1 U13 ( .A1(n1), .A2(IN1[12]), .ZN(n15) );
  NAND2_X1 U14 ( .A1(n9), .A2(n15), .ZN(Y[12]) );
  NAND2_X1 U15 ( .A1(n1), .A2(IN1[13]), .ZN(n16) );
  NAND2_X1 U16 ( .A1(n9), .A2(n16), .ZN(Y[13]) );
  NAND2_X1 U17 ( .A1(n1), .A2(IN1[14]), .ZN(n17) );
  NAND2_X1 U18 ( .A1(n9), .A2(n17), .ZN(Y[14]) );
  NAND2_X1 U19 ( .A1(n1), .A2(IN1[15]), .ZN(n18) );
  NAND2_X1 U20 ( .A1(n9), .A2(n18), .ZN(Y[15]) );
  NAND2_X1 U21 ( .A1(n1), .A2(IN1[16]), .ZN(n19) );
  NAND2_X1 U22 ( .A1(n9), .A2(n19), .ZN(Y[16]) );
  NAND2_X1 U23 ( .A1(n1), .A2(IN1[17]), .ZN(n20) );
  NAND2_X1 U24 ( .A1(n9), .A2(n20), .ZN(Y[17]) );
  NAND2_X1 U25 ( .A1(n1), .A2(IN1[18]), .ZN(n21) );
  NAND2_X1 U26 ( .A1(n9), .A2(n21), .ZN(Y[18]) );
  NAND2_X1 U27 ( .A1(n1), .A2(IN1[19]), .ZN(n22) );
  NAND2_X1 U28 ( .A1(n9), .A2(n22), .ZN(Y[19]) );
  NAND2_X1 U29 ( .A1(n1), .A2(IN1[1]), .ZN(n23) );
  NAND2_X1 U30 ( .A1(n1), .A2(IN1[20]), .ZN(n24) );
  NAND2_X1 U31 ( .A1(n9), .A2(n24), .ZN(Y[20]) );
  NAND2_X1 U32 ( .A1(n1), .A2(IN1[21]), .ZN(n25) );
  NAND2_X1 U33 ( .A1(n9), .A2(n25), .ZN(Y[21]) );
  NAND2_X1 U34 ( .A1(n1), .A2(IN1[22]), .ZN(n26) );
  NAND2_X1 U35 ( .A1(n9), .A2(n26), .ZN(Y[22]) );
  NAND2_X1 U36 ( .A1(n1), .A2(IN1[23]), .ZN(n27) );
  NAND2_X1 U37 ( .A1(n9), .A2(n27), .ZN(Y[23]) );
  NAND2_X1 U38 ( .A1(n1), .A2(IN1[24]), .ZN(n28) );
  NAND2_X1 U39 ( .A1(n9), .A2(n28), .ZN(Y[24]) );
  NAND2_X1 U40 ( .A1(n1), .A2(IN1[25]), .ZN(n29) );
  NAND2_X1 U41 ( .A1(n9), .A2(n29), .ZN(Y[25]) );
  NAND2_X1 U42 ( .A1(n1), .A2(IN1[26]), .ZN(n30) );
  NAND2_X1 U43 ( .A1(n10), .A2(n30), .ZN(Y[26]) );
  NAND2_X1 U44 ( .A1(n1), .A2(IN1[27]), .ZN(n31) );
  NAND2_X1 U45 ( .A1(n9), .A2(n31), .ZN(Y[27]) );
  NAND2_X1 U46 ( .A1(n1), .A2(IN1[28]), .ZN(n32) );
  NAND2_X1 U47 ( .A1(n9), .A2(n32), .ZN(Y[28]) );
  NAND2_X1 U48 ( .A1(n1), .A2(IN1[29]), .ZN(n33) );
  NAND2_X1 U49 ( .A1(n9), .A2(n33), .ZN(Y[29]) );
  NAND2_X1 U50 ( .A1(n1), .A2(IN1[2]), .ZN(n34) );
  NAND2_X1 U51 ( .A1(n10), .A2(n34), .ZN(Y[2]) );
  NAND2_X1 U52 ( .A1(n1), .A2(IN1[30]), .ZN(n35) );
  NAND2_X1 U53 ( .A1(n10), .A2(n35), .ZN(Y[30]) );
  NAND2_X1 U54 ( .A1(n1), .A2(IN1[3]), .ZN(n36) );
  NAND2_X1 U55 ( .A1(n10), .A2(n36), .ZN(Y[3]) );
  NAND2_X1 U56 ( .A1(n1), .A2(IN1[4]), .ZN(n37) );
  NAND2_X1 U57 ( .A1(n10), .A2(n37), .ZN(Y[4]) );
  NAND2_X1 U58 ( .A1(n1), .A2(IN1[5]), .ZN(n38) );
  NAND2_X1 U59 ( .A1(n10), .A2(n38), .ZN(Y[5]) );
  NAND2_X1 U60 ( .A1(n1), .A2(IN1[6]), .ZN(n39) );
  NAND2_X1 U61 ( .A1(n10), .A2(n39), .ZN(Y[6]) );
  NAND2_X1 U62 ( .A1(n1), .A2(IN1[7]), .ZN(n40) );
  NAND2_X1 U63 ( .A1(n10), .A2(n40), .ZN(Y[7]) );
  NAND2_X1 U64 ( .A1(n1), .A2(IN1[8]), .ZN(n41) );
  NAND2_X1 U65 ( .A1(n10), .A2(n41), .ZN(Y[8]) );
  NAND2_X1 U66 ( .A1(n1), .A2(IN1[9]), .ZN(n42) );
  NAND2_X1 U67 ( .A1(n10), .A2(n42), .ZN(Y[9]) );
endmodule


module MUX_2to1_N4_0 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  AND2_X1 U1 ( .A1(SEL), .A2(IN1[0]), .ZN(Y[0]) );
  AND2_X1 U2 ( .A1(SEL), .A2(IN1[1]), .ZN(Y[1]) );
  AND2_X1 U3 ( .A1(SEL), .A2(IN1[2]), .ZN(Y[2]) );
  AND2_X1 U4 ( .A1(SEL), .A2(IN1[3]), .ZN(Y[3]) );
endmodule


module MUX_2to1_N8 ( IN0, IN1, SEL, Y );
  input [7:0] IN0;
  input [7:0] IN1;
  output [7:0] Y;
  input SEL;


  AND2_X1 U1 ( .A1(SEL), .A2(IN1[0]), .ZN(Y[0]) );
  AND2_X1 U2 ( .A1(SEL), .A2(IN1[1]), .ZN(Y[1]) );
  AND2_X1 U3 ( .A1(SEL), .A2(IN1[2]), .ZN(Y[2]) );
  AND2_X1 U4 ( .A1(SEL), .A2(IN1[3]), .ZN(Y[3]) );
  AND2_X1 U5 ( .A1(SEL), .A2(IN1[4]), .ZN(Y[4]) );
  AND2_X1 U6 ( .A1(SEL), .A2(IN1[5]), .ZN(Y[5]) );
  AND2_X1 U7 ( .A1(SEL), .A2(IN1[6]), .ZN(Y[6]) );
  AND2_X1 U8 ( .A1(SEL), .A2(IN1[7]), .ZN(Y[7]) );
endmodule


module MUX_2to1_N12 ( IN0, IN1, SEL, Y );
  input [11:0] IN0;
  input [11:0] IN1;
  output [11:0] Y;
  input SEL;


  AND2_X1 U1 ( .A1(SEL), .A2(IN1[0]), .ZN(Y[0]) );
  AND2_X1 U2 ( .A1(SEL), .A2(IN1[1]), .ZN(Y[1]) );
  AND2_X1 U3 ( .A1(SEL), .A2(IN1[2]), .ZN(Y[2]) );
  AND2_X1 U4 ( .A1(SEL), .A2(IN1[3]), .ZN(Y[3]) );
  AND2_X1 U5 ( .A1(SEL), .A2(IN1[4]), .ZN(Y[4]) );
  AND2_X1 U6 ( .A1(SEL), .A2(IN1[5]), .ZN(Y[5]) );
  AND2_X1 U7 ( .A1(SEL), .A2(IN1[6]), .ZN(Y[6]) );
  AND2_X1 U8 ( .A1(SEL), .A2(IN1[7]), .ZN(Y[7]) );
  AND2_X1 U9 ( .A1(SEL), .A2(IN1[8]), .ZN(Y[8]) );
  AND2_X1 U10 ( .A1(SEL), .A2(IN1[9]), .ZN(Y[9]) );
  AND2_X1 U11 ( .A1(SEL), .A2(IN1[10]), .ZN(Y[10]) );
  AND2_X1 U12 ( .A1(SEL), .A2(IN1[11]), .ZN(Y[11]) );
endmodule


module MUX_2to1_N16 ( IN0, IN1, SEL, Y );
  input [15:0] IN0;
  input [15:0] IN1;
  output [15:0] Y;
  input SEL;


  AND2_X1 U1 ( .A1(SEL), .A2(IN1[0]), .ZN(Y[0]) );
  AND2_X1 U2 ( .A1(SEL), .A2(IN1[1]), .ZN(Y[1]) );
  AND2_X1 U3 ( .A1(SEL), .A2(IN1[2]), .ZN(Y[2]) );
  AND2_X1 U4 ( .A1(SEL), .A2(IN1[3]), .ZN(Y[3]) );
  AND2_X1 U5 ( .A1(SEL), .A2(IN1[4]), .ZN(Y[4]) );
  AND2_X1 U6 ( .A1(SEL), .A2(IN1[5]), .ZN(Y[5]) );
  AND2_X1 U7 ( .A1(SEL), .A2(IN1[6]), .ZN(Y[6]) );
  AND2_X1 U8 ( .A1(SEL), .A2(IN1[7]), .ZN(Y[7]) );
  AND2_X1 U9 ( .A1(SEL), .A2(IN1[8]), .ZN(Y[8]) );
  AND2_X1 U10 ( .A1(SEL), .A2(IN1[9]), .ZN(Y[9]) );
  AND2_X1 U11 ( .A1(SEL), .A2(IN1[10]), .ZN(Y[10]) );
  AND2_X1 U12 ( .A1(SEL), .A2(IN1[11]), .ZN(Y[11]) );
  AND2_X1 U13 ( .A1(SEL), .A2(IN1[12]), .ZN(Y[12]) );
  AND2_X1 U14 ( .A1(SEL), .A2(IN1[13]), .ZN(Y[13]) );
  AND2_X1 U15 ( .A1(SEL), .A2(IN1[14]), .ZN(Y[14]) );
  AND2_X1 U16 ( .A1(SEL), .A2(IN1[15]), .ZN(Y[15]) );
endmodule


module MUX_2to1_N20 ( IN0, IN1, SEL, Y );
  input [19:0] IN0;
  input [19:0] IN1;
  output [19:0] Y;
  input SEL;


  AND2_X1 U1 ( .A1(SEL), .A2(IN1[0]), .ZN(Y[0]) );
  AND2_X1 U2 ( .A1(SEL), .A2(IN1[1]), .ZN(Y[1]) );
  AND2_X1 U3 ( .A1(SEL), .A2(IN1[2]), .ZN(Y[2]) );
  AND2_X1 U4 ( .A1(SEL), .A2(IN1[3]), .ZN(Y[3]) );
  AND2_X1 U5 ( .A1(SEL), .A2(IN1[4]), .ZN(Y[4]) );
  AND2_X1 U6 ( .A1(SEL), .A2(IN1[5]), .ZN(Y[5]) );
  AND2_X1 U7 ( .A1(SEL), .A2(IN1[6]), .ZN(Y[6]) );
  AND2_X1 U8 ( .A1(SEL), .A2(IN1[7]), .ZN(Y[7]) );
  AND2_X1 U9 ( .A1(SEL), .A2(IN1[8]), .ZN(Y[8]) );
  AND2_X1 U10 ( .A1(SEL), .A2(IN1[9]), .ZN(Y[9]) );
  AND2_X1 U11 ( .A1(SEL), .A2(IN1[10]), .ZN(Y[10]) );
  AND2_X1 U12 ( .A1(SEL), .A2(IN1[11]), .ZN(Y[11]) );
  AND2_X1 U13 ( .A1(SEL), .A2(IN1[12]), .ZN(Y[12]) );
  AND2_X1 U14 ( .A1(SEL), .A2(IN1[13]), .ZN(Y[13]) );
  AND2_X1 U15 ( .A1(SEL), .A2(IN1[14]), .ZN(Y[14]) );
  AND2_X1 U16 ( .A1(SEL), .A2(IN1[15]), .ZN(Y[15]) );
  AND2_X1 U17 ( .A1(SEL), .A2(IN1[16]), .ZN(Y[16]) );
  AND2_X1 U18 ( .A1(SEL), .A2(IN1[17]), .ZN(Y[17]) );
  AND2_X1 U19 ( .A1(SEL), .A2(IN1[18]), .ZN(Y[18]) );
  AND2_X1 U20 ( .A1(SEL), .A2(IN1[19]), .ZN(Y[19]) );
endmodule


module MUX_2to1_N24 ( IN0, IN1, SEL, Y );
  input [23:0] IN0;
  input [23:0] IN1;
  output [23:0] Y;
  input SEL;
  wire   n1;

  BUF_X2 U1 ( .A(SEL), .Z(n1) );
  AND2_X1 U2 ( .A1(n1), .A2(IN1[0]), .ZN(Y[0]) );
  AND2_X1 U3 ( .A1(SEL), .A2(IN1[1]), .ZN(Y[1]) );
  AND2_X1 U4 ( .A1(n1), .A2(IN1[2]), .ZN(Y[2]) );
  AND2_X1 U5 ( .A1(n1), .A2(IN1[3]), .ZN(Y[3]) );
  AND2_X1 U6 ( .A1(n1), .A2(IN1[4]), .ZN(Y[4]) );
  AND2_X1 U7 ( .A1(n1), .A2(IN1[5]), .ZN(Y[5]) );
  AND2_X1 U8 ( .A1(n1), .A2(IN1[6]), .ZN(Y[6]) );
  AND2_X1 U9 ( .A1(n1), .A2(IN1[7]), .ZN(Y[7]) );
  AND2_X1 U10 ( .A1(n1), .A2(IN1[8]), .ZN(Y[8]) );
  AND2_X1 U11 ( .A1(n1), .A2(IN1[9]), .ZN(Y[9]) );
  AND2_X1 U12 ( .A1(n1), .A2(IN1[10]), .ZN(Y[10]) );
  AND2_X1 U13 ( .A1(n1), .A2(IN1[11]), .ZN(Y[11]) );
  AND2_X1 U14 ( .A1(n1), .A2(IN1[12]), .ZN(Y[12]) );
  AND2_X1 U15 ( .A1(n1), .A2(IN1[13]), .ZN(Y[13]) );
  AND2_X1 U16 ( .A1(SEL), .A2(IN1[14]), .ZN(Y[14]) );
  AND2_X1 U17 ( .A1(n1), .A2(IN1[15]), .ZN(Y[15]) );
  AND2_X1 U18 ( .A1(n1), .A2(IN1[16]), .ZN(Y[16]) );
  AND2_X1 U19 ( .A1(n1), .A2(IN1[17]), .ZN(Y[17]) );
  AND2_X1 U20 ( .A1(SEL), .A2(IN1[18]), .ZN(Y[18]) );
  AND2_X1 U21 ( .A1(n1), .A2(IN1[19]), .ZN(Y[19]) );
  AND2_X1 U22 ( .A1(SEL), .A2(IN1[20]), .ZN(Y[20]) );
  AND2_X1 U23 ( .A1(SEL), .A2(IN1[21]), .ZN(Y[21]) );
  AND2_X1 U24 ( .A1(n1), .A2(IN1[22]), .ZN(Y[22]) );
  AND2_X1 U25 ( .A1(n1), .A2(IN1[23]), .ZN(Y[23]) );
endmodule


module MUX_2to1_N28 ( IN0, IN1, SEL, Y );
  input [27:0] IN0;
  input [27:0] IN1;
  output [27:0] Y;
  input SEL;
  wire   n1;

  AND2_X1 U1 ( .A1(IN1[1]), .A2(SEL), .ZN(Y[1]) );
  BUF_X1 U2 ( .A(SEL), .Z(n1) );
  AND2_X1 U3 ( .A1(SEL), .A2(IN1[0]), .ZN(Y[0]) );
  AND2_X1 U4 ( .A1(SEL), .A2(IN1[2]), .ZN(Y[2]) );
  AND2_X1 U5 ( .A1(SEL), .A2(IN1[3]), .ZN(Y[3]) );
  AND2_X1 U6 ( .A1(SEL), .A2(IN1[4]), .ZN(Y[4]) );
  AND2_X1 U7 ( .A1(SEL), .A2(IN1[5]), .ZN(Y[5]) );
  AND2_X1 U8 ( .A1(SEL), .A2(IN1[6]), .ZN(Y[6]) );
  AND2_X1 U9 ( .A1(SEL), .A2(IN1[7]), .ZN(Y[7]) );
  AND2_X1 U10 ( .A1(n1), .A2(IN1[8]), .ZN(Y[8]) );
  AND2_X1 U11 ( .A1(n1), .A2(IN1[9]), .ZN(Y[9]) );
  AND2_X1 U12 ( .A1(n1), .A2(IN1[10]), .ZN(Y[10]) );
  AND2_X1 U13 ( .A1(n1), .A2(IN1[11]), .ZN(Y[11]) );
  AND2_X1 U14 ( .A1(n1), .A2(IN1[12]), .ZN(Y[12]) );
  AND2_X1 U15 ( .A1(n1), .A2(IN1[13]), .ZN(Y[13]) );
  AND2_X1 U16 ( .A1(n1), .A2(IN1[14]), .ZN(Y[14]) );
  AND2_X1 U17 ( .A1(n1), .A2(IN1[15]), .ZN(Y[15]) );
  AND2_X1 U18 ( .A1(n1), .A2(IN1[16]), .ZN(Y[16]) );
  AND2_X1 U19 ( .A1(n1), .A2(IN1[17]), .ZN(Y[17]) );
  AND2_X1 U20 ( .A1(n1), .A2(IN1[18]), .ZN(Y[18]) );
  AND2_X1 U21 ( .A1(SEL), .A2(IN1[19]), .ZN(Y[19]) );
  AND2_X1 U22 ( .A1(n1), .A2(IN1[20]), .ZN(Y[20]) );
  AND2_X1 U23 ( .A1(SEL), .A2(IN1[21]), .ZN(Y[21]) );
  AND2_X1 U24 ( .A1(SEL), .A2(IN1[22]), .ZN(Y[22]) );
  AND2_X1 U25 ( .A1(SEL), .A2(IN1[23]), .ZN(Y[23]) );
  AND2_X1 U26 ( .A1(SEL), .A2(IN1[24]), .ZN(Y[24]) );
  AND2_X1 U27 ( .A1(SEL), .A2(IN1[25]), .ZN(Y[25]) );
  AND2_X1 U28 ( .A1(SEL), .A2(IN1[26]), .ZN(Y[26]) );
  AND2_X1 U29 ( .A1(SEL), .A2(IN1[27]), .ZN(Y[27]) );
endmodule


module MUX_2to1_N32_2 ( IN0, IN1, SEL, Y );
  input [31:0] IN0;
  input [31:0] IN1;
  output [31:0] Y;
  input SEL;


  AND2_X1 U1 ( .A1(SEL), .A2(IN1[0]), .ZN(Y[0]) );
  AND2_X1 U2 ( .A1(SEL), .A2(IN1[1]), .ZN(Y[1]) );
  AND2_X1 U3 ( .A1(SEL), .A2(IN1[2]), .ZN(Y[2]) );
  AND2_X1 U4 ( .A1(SEL), .A2(IN1[3]), .ZN(Y[3]) );
  AND2_X1 U5 ( .A1(SEL), .A2(IN1[4]), .ZN(Y[4]) );
  AND2_X1 U6 ( .A1(SEL), .A2(IN1[5]), .ZN(Y[5]) );
  AND2_X1 U7 ( .A1(SEL), .A2(IN1[6]), .ZN(Y[6]) );
  AND2_X1 U8 ( .A1(SEL), .A2(IN1[7]), .ZN(Y[7]) );
  AND2_X1 U9 ( .A1(SEL), .A2(IN1[8]), .ZN(Y[8]) );
  AND2_X1 U10 ( .A1(SEL), .A2(IN1[9]), .ZN(Y[9]) );
  AND2_X1 U11 ( .A1(SEL), .A2(IN1[10]), .ZN(Y[10]) );
  AND2_X1 U12 ( .A1(SEL), .A2(IN1[11]), .ZN(Y[11]) );
  AND2_X1 U13 ( .A1(SEL), .A2(IN1[12]), .ZN(Y[12]) );
  AND2_X1 U14 ( .A1(SEL), .A2(IN1[13]), .ZN(Y[13]) );
  AND2_X1 U15 ( .A1(SEL), .A2(IN1[14]), .ZN(Y[14]) );
  AND2_X1 U16 ( .A1(SEL), .A2(IN1[15]), .ZN(Y[15]) );
  AND2_X1 U17 ( .A1(SEL), .A2(IN1[16]), .ZN(Y[16]) );
  AND2_X1 U18 ( .A1(SEL), .A2(IN1[17]), .ZN(Y[17]) );
  AND2_X1 U19 ( .A1(SEL), .A2(IN1[18]), .ZN(Y[18]) );
  AND2_X1 U20 ( .A1(SEL), .A2(IN1[19]), .ZN(Y[19]) );
  AND2_X1 U21 ( .A1(SEL), .A2(IN1[20]), .ZN(Y[20]) );
  AND2_X1 U22 ( .A1(SEL), .A2(IN1[21]), .ZN(Y[21]) );
  AND2_X1 U23 ( .A1(SEL), .A2(IN1[22]), .ZN(Y[22]) );
  AND2_X1 U24 ( .A1(SEL), .A2(IN1[23]), .ZN(Y[23]) );
  AND2_X1 U25 ( .A1(SEL), .A2(IN1[24]), .ZN(Y[24]) );
  AND2_X1 U26 ( .A1(SEL), .A2(IN1[25]), .ZN(Y[25]) );
  AND2_X1 U27 ( .A1(SEL), .A2(IN1[26]), .ZN(Y[26]) );
  AND2_X1 U28 ( .A1(SEL), .A2(IN1[27]), .ZN(Y[27]) );
  AND2_X1 U29 ( .A1(SEL), .A2(IN1[28]), .ZN(Y[28]) );
  AND2_X1 U30 ( .A1(SEL), .A2(IN1[29]), .ZN(Y[29]) );
  AND2_X1 U31 ( .A1(SEL), .A2(IN1[30]), .ZN(Y[30]) );
  AND2_X1 U32 ( .A1(SEL), .A2(IN1[31]), .ZN(Y[31]) );
endmodule


module MUX_2to1_N36_0 ( IN0, IN1, SEL, Y );
  input [35:0] IN0;
  input [35:0] IN1;
  output [35:0] Y;
  input SEL;
  wire   n8, n9, n10;

  OAI21_X1 U1 ( .B1(n10), .B2(n9), .A(n8), .ZN(Y[9]) );
  NAND2_X1 U2 ( .A1(n10), .A2(IN0[13]), .ZN(n8) );
  INV_X1 U3 ( .A(IN1[5]), .ZN(n9) );
  BUF_X1 U4 ( .A(SEL), .Z(n10) );
  MUX2_X1 U5 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U6 ( .A(IN0[10]), .B(IN1[10]), .S(SEL), .Z(Y[10]) );
  MUX2_X1 U7 ( .A(IN0[11]), .B(IN1[11]), .S(SEL), .Z(Y[11]) );
  MUX2_X1 U8 ( .A(IN0[12]), .B(IN1[12]), .S(SEL), .Z(Y[12]) );
  MUX2_X1 U9 ( .A(IN0[13]), .B(IN1[13]), .S(SEL), .Z(Y[13]) );
  MUX2_X1 U10 ( .A(IN1[10]), .B(IN1[14]), .S(SEL), .Z(Y[14]) );
  MUX2_X1 U11 ( .A(IN1[11]), .B(IN1[15]), .S(SEL), .Z(Y[15]) );
  MUX2_X1 U12 ( .A(IN1[12]), .B(IN1[16]), .S(SEL), .Z(Y[16]) );
  MUX2_X1 U13 ( .A(IN1[13]), .B(IN1[17]), .S(SEL), .Z(Y[17]) );
  MUX2_X1 U14 ( .A(IN1[14]), .B(IN1[18]), .S(SEL), .Z(Y[18]) );
  MUX2_X1 U15 ( .A(IN1[15]), .B(IN1[19]), .S(SEL), .Z(Y[19]) );
  MUX2_X1 U16 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U17 ( .A(IN1[16]), .B(IN1[20]), .S(SEL), .Z(Y[20]) );
  MUX2_X1 U18 ( .A(IN1[17]), .B(IN1[21]), .S(SEL), .Z(Y[21]) );
  MUX2_X1 U19 ( .A(IN1[18]), .B(IN1[22]), .S(SEL), .Z(Y[22]) );
  MUX2_X1 U20 ( .A(IN1[19]), .B(IN1[23]), .S(SEL), .Z(Y[23]) );
  MUX2_X1 U21 ( .A(IN1[20]), .B(IN1[24]), .S(SEL), .Z(Y[24]) );
  MUX2_X1 U22 ( .A(IN1[21]), .B(IN1[25]), .S(SEL), .Z(Y[25]) );
  MUX2_X1 U23 ( .A(IN1[22]), .B(IN1[26]), .S(SEL), .Z(Y[26]) );
  MUX2_X1 U24 ( .A(IN1[23]), .B(IN1[27]), .S(SEL), .Z(Y[27]) );
  MUX2_X1 U25 ( .A(IN1[24]), .B(IN1[28]), .S(SEL), .Z(Y[28]) );
  MUX2_X1 U26 ( .A(IN1[25]), .B(IN1[29]), .S(SEL), .Z(Y[29]) );
  MUX2_X1 U27 ( .A(IN0[2]), .B(IN1[2]), .S(n10), .Z(Y[2]) );
  MUX2_X1 U28 ( .A(IN1[26]), .B(IN1[30]), .S(n10), .Z(Y[30]) );
  MUX2_X1 U29 ( .A(IN1[27]), .B(IN1[31]), .S(n10), .Z(Y[31]) );
  MUX2_X1 U30 ( .A(IN1[28]), .B(IN1[32]), .S(n10), .Z(Y[32]) );
  MUX2_X1 U31 ( .A(IN1[29]), .B(IN1[33]), .S(n10), .Z(Y[33]) );
  MUX2_X1 U32 ( .A(IN1[30]), .B(IN1[34]), .S(n10), .Z(Y[34]) );
  MUX2_X1 U33 ( .A(IN1[31]), .B(IN1[35]), .S(n10), .Z(Y[35]) );
  MUX2_X1 U34 ( .A(IN0[3]), .B(IN1[3]), .S(n10), .Z(Y[3]) );
  MUX2_X1 U35 ( .A(IN1[0]), .B(IN1[4]), .S(n10), .Z(Y[4]) );
  MUX2_X1 U36 ( .A(IN1[1]), .B(IN1[5]), .S(n10), .Z(Y[5]) );
  MUX2_X1 U37 ( .A(IN1[2]), .B(IN0[10]), .S(n10), .Z(Y[6]) );
  MUX2_X1 U38 ( .A(IN1[3]), .B(IN0[11]), .S(n10), .Z(Y[7]) );
  MUX2_X1 U39 ( .A(IN1[4]), .B(IN0[12]), .S(n10), .Z(Y[8]) );
endmodule


module MUX_2to1_N36_7 ( IN0, IN1, SEL, Y );
  input [35:0] IN0;
  input [35:0] IN1;
  output [35:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(IN0[10]), .B(IN1[10]), .S(SEL), .Z(Y[10]) );
  MUX2_X1 U3 ( .A(IN0[11]), .B(IN1[11]), .S(SEL), .Z(Y[11]) );
  MUX2_X1 U4 ( .A(IN1[0]), .B(IN1[12]), .S(SEL), .Z(Y[12]) );
  MUX2_X1 U5 ( .A(IN0[13]), .B(IN1[13]), .S(SEL), .Z(Y[13]) );
  MUX2_X1 U6 ( .A(IN0[14]), .B(IN1[14]), .S(SEL), .Z(Y[14]) );
  MUX2_X1 U7 ( .A(IN0[15]), .B(IN1[15]), .S(SEL), .Z(Y[15]) );
  MUX2_X1 U8 ( .A(IN0[16]), .B(IN1[16]), .S(SEL), .Z(Y[16]) );
  MUX2_X1 U9 ( .A(IN0[17]), .B(IN1[17]), .S(SEL), .Z(Y[17]) );
  MUX2_X1 U10 ( .A(IN0[18]), .B(IN1[18]), .S(SEL), .Z(Y[18]) );
  MUX2_X1 U11 ( .A(IN0[19]), .B(IN1[19]), .S(SEL), .Z(Y[19]) );
  MUX2_X1 U12 ( .A(IN0[1]), .B(IN0[13]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U13 ( .A(IN0[20]), .B(IN1[20]), .S(SEL), .Z(Y[20]) );
  MUX2_X1 U14 ( .A(IN0[21]), .B(IN1[21]), .S(SEL), .Z(Y[21]) );
  MUX2_X1 U15 ( .A(IN1[10]), .B(IN1[22]), .S(SEL), .Z(Y[22]) );
  MUX2_X1 U16 ( .A(IN1[11]), .B(IN1[23]), .S(SEL), .Z(Y[23]) );
  MUX2_X1 U17 ( .A(IN1[12]), .B(IN1[24]), .S(SEL), .Z(Y[24]) );
  MUX2_X1 U18 ( .A(IN1[13]), .B(IN1[25]), .S(SEL), .Z(Y[25]) );
  MUX2_X1 U19 ( .A(IN1[14]), .B(IN1[26]), .S(SEL), .Z(Y[26]) );
  MUX2_X1 U20 ( .A(IN1[15]), .B(IN1[27]), .S(SEL), .Z(Y[27]) );
  MUX2_X1 U21 ( .A(IN1[16]), .B(IN1[28]), .S(SEL), .Z(Y[28]) );
  MUX2_X1 U22 ( .A(IN1[17]), .B(IN1[29]), .S(SEL), .Z(Y[29]) );
  MUX2_X1 U23 ( .A(IN0[2]), .B(IN0[14]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U24 ( .A(IN1[18]), .B(IN1[30]), .S(SEL), .Z(Y[30]) );
  MUX2_X1 U25 ( .A(IN1[19]), .B(IN1[31]), .S(SEL), .Z(Y[31]) );
  MUX2_X1 U26 ( .A(IN1[20]), .B(IN1[32]), .S(SEL), .Z(Y[32]) );
  MUX2_X1 U27 ( .A(IN1[21]), .B(IN1[33]), .S(SEL), .Z(Y[33]) );
  MUX2_X1 U28 ( .A(IN1[22]), .B(IN1[34]), .S(SEL), .Z(Y[34]) );
  MUX2_X1 U29 ( .A(IN1[23]), .B(IN1[35]), .S(SEL), .Z(Y[35]) );
  MUX2_X1 U30 ( .A(IN0[3]), .B(IN0[15]), .S(SEL), .Z(Y[3]) );
  MUX2_X1 U31 ( .A(IN0[4]), .B(IN0[16]), .S(SEL), .Z(Y[4]) );
  MUX2_X1 U32 ( .A(IN0[5]), .B(IN0[17]), .S(SEL), .Z(Y[5]) );
  MUX2_X1 U33 ( .A(IN0[6]), .B(IN0[18]), .S(SEL), .Z(Y[6]) );
  MUX2_X1 U34 ( .A(IN0[7]), .B(IN0[19]), .S(SEL), .Z(Y[7]) );
  MUX2_X1 U35 ( .A(IN0[8]), .B(IN0[20]), .S(SEL), .Z(Y[8]) );
  MUX2_X1 U36 ( .A(IN0[9]), .B(IN0[21]), .S(SEL), .Z(Y[9]) );
endmodule


module MUX_2to1_N36_6 ( IN0, IN1, SEL, Y );
  input [35:0] IN0;
  input [35:0] IN1;
  output [35:0] Y;
  input SEL;
  wire   n8, n9, n10, n11;

  BUF_X2 U1 ( .A(SEL), .Z(n10) );
  NAND2_X1 U2 ( .A1(n11), .A2(IN0[29]), .ZN(n8) );
  OAI21_X1 U3 ( .B1(n10), .B2(n9), .A(n8), .ZN(Y[9]) );
  INV_X1 U4 ( .A(IN0[9]), .ZN(n9) );
  BUF_X1 U5 ( .A(SEL), .Z(n11) );
  MUX2_X1 U6 ( .A(IN0[0]), .B(IN1[0]), .S(n11), .Z(Y[0]) );
  MUX2_X1 U7 ( .A(IN0[10]), .B(IN1[10]), .S(SEL), .Z(Y[10]) );
  MUX2_X1 U8 ( .A(IN0[11]), .B(IN1[11]), .S(SEL), .Z(Y[11]) );
  MUX2_X1 U9 ( .A(IN0[12]), .B(IN1[12]), .S(SEL), .Z(Y[12]) );
  MUX2_X1 U10 ( .A(IN0[13]), .B(IN1[13]), .S(SEL), .Z(Y[13]) );
  MUX2_X1 U11 ( .A(IN0[14]), .B(IN1[14]), .S(SEL), .Z(Y[14]) );
  MUX2_X1 U12 ( .A(IN0[15]), .B(IN1[15]), .S(SEL), .Z(Y[15]) );
  MUX2_X1 U13 ( .A(IN0[16]), .B(IN1[16]), .S(SEL), .Z(Y[16]) );
  MUX2_X1 U14 ( .A(IN0[17]), .B(IN1[17]), .S(n10), .Z(Y[17]) );
  MUX2_X1 U15 ( .A(IN0[18]), .B(IN1[18]), .S(n10), .Z(Y[18]) );
  MUX2_X1 U16 ( .A(IN0[19]), .B(IN1[19]), .S(n10), .Z(Y[19]) );
  MUX2_X1 U17 ( .A(IN0[1]), .B(IN1[1]), .S(n11), .Z(Y[1]) );
  MUX2_X1 U18 ( .A(IN1[0]), .B(IN1[20]), .S(n10), .Z(Y[20]) );
  MUX2_X1 U19 ( .A(IN1[1]), .B(IN1[21]), .S(SEL), .Z(Y[21]) );
  MUX2_X1 U20 ( .A(IN0[22]), .B(IN1[22]), .S(n10), .Z(Y[22]) );
  MUX2_X1 U21 ( .A(IN0[23]), .B(IN1[23]), .S(n10), .Z(Y[23]) );
  MUX2_X1 U22 ( .A(IN0[24]), .B(IN1[24]), .S(n11), .Z(Y[24]) );
  MUX2_X1 U23 ( .A(IN0[25]), .B(IN1[25]), .S(n10), .Z(Y[25]) );
  MUX2_X1 U24 ( .A(IN0[26]), .B(IN1[26]), .S(n11), .Z(Y[26]) );
  MUX2_X1 U25 ( .A(IN0[27]), .B(IN1[27]), .S(n10), .Z(Y[27]) );
  MUX2_X1 U26 ( .A(IN0[28]), .B(IN1[28]), .S(n11), .Z(Y[28]) );
  MUX2_X1 U27 ( .A(IN0[29]), .B(IN1[29]), .S(n10), .Z(Y[29]) );
  MUX2_X1 U28 ( .A(IN0[2]), .B(IN0[22]), .S(n11), .Z(Y[2]) );
  MUX2_X1 U29 ( .A(IN1[10]), .B(IN1[30]), .S(n11), .Z(Y[30]) );
  MUX2_X1 U30 ( .A(IN1[11]), .B(IN1[31]), .S(n10), .Z(Y[31]) );
  MUX2_X1 U31 ( .A(IN1[12]), .B(IN1[32]), .S(n11), .Z(Y[32]) );
  MUX2_X1 U32 ( .A(IN1[13]), .B(IN1[33]), .S(n11), .Z(Y[33]) );
  MUX2_X1 U33 ( .A(IN1[14]), .B(IN1[34]), .S(n11), .Z(Y[34]) );
  MUX2_X1 U34 ( .A(IN1[15]), .B(IN1[35]), .S(n11), .Z(Y[35]) );
  MUX2_X1 U35 ( .A(IN0[3]), .B(IN0[23]), .S(n11), .Z(Y[3]) );
  MUX2_X1 U36 ( .A(IN0[4]), .B(IN0[24]), .S(n11), .Z(Y[4]) );
  MUX2_X1 U37 ( .A(IN0[5]), .B(IN0[25]), .S(n11), .Z(Y[5]) );
  MUX2_X1 U38 ( .A(IN0[6]), .B(IN0[26]), .S(n11), .Z(Y[6]) );
  MUX2_X1 U39 ( .A(IN0[7]), .B(IN0[27]), .S(n10), .Z(Y[7]) );
  MUX2_X1 U40 ( .A(IN0[8]), .B(IN0[28]), .S(n10), .Z(Y[8]) );
endmodule


module MUX_2to1_N36_5 ( IN0, IN1, SEL, Y );
  input [35:0] IN0;
  input [35:0] IN1;
  output [35:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(IN0[10]), .B(IN1[10]), .S(SEL), .Z(Y[10]) );
  MUX2_X1 U3 ( .A(IN0[11]), .B(IN1[11]), .S(SEL), .Z(Y[11]) );
  MUX2_X1 U4 ( .A(IN0[12]), .B(IN1[12]), .S(SEL), .Z(Y[12]) );
  MUX2_X1 U5 ( .A(IN0[13]), .B(IN1[13]), .S(SEL), .Z(Y[13]) );
  MUX2_X1 U6 ( .A(IN0[14]), .B(IN1[14]), .S(SEL), .Z(Y[14]) );
  MUX2_X1 U7 ( .A(IN0[15]), .B(IN1[15]), .S(SEL), .Z(Y[15]) );
  MUX2_X1 U8 ( .A(IN0[16]), .B(IN1[16]), .S(SEL), .Z(Y[16]) );
  MUX2_X1 U9 ( .A(IN0[17]), .B(IN1[17]), .S(SEL), .Z(Y[17]) );
  MUX2_X1 U10 ( .A(IN0[18]), .B(IN1[18]), .S(SEL), .Z(Y[18]) );
  MUX2_X1 U11 ( .A(IN0[19]), .B(IN1[19]), .S(SEL), .Z(Y[19]) );
  MUX2_X1 U12 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U13 ( .A(IN0[20]), .B(IN1[20]), .S(SEL), .Z(Y[20]) );
  MUX2_X1 U14 ( .A(IN0[21]), .B(IN1[21]), .S(SEL), .Z(Y[21]) );
  MUX2_X1 U15 ( .A(IN0[22]), .B(IN1[22]), .S(SEL), .Z(Y[22]) );
  MUX2_X1 U16 ( .A(IN0[23]), .B(IN1[23]), .S(SEL), .Z(Y[23]) );
  MUX2_X1 U17 ( .A(IN0[24]), .B(IN1[24]), .S(SEL), .Z(Y[24]) );
  MUX2_X1 U18 ( .A(IN0[25]), .B(IN1[25]), .S(SEL), .Z(Y[25]) );
  MUX2_X1 U19 ( .A(IN0[26]), .B(IN1[26]), .S(SEL), .Z(Y[26]) );
  MUX2_X1 U20 ( .A(IN0[27]), .B(IN1[27]), .S(SEL), .Z(Y[27]) );
  MUX2_X1 U21 ( .A(IN1[0]), .B(IN1[28]), .S(SEL), .Z(Y[28]) );
  MUX2_X1 U22 ( .A(IN1[1]), .B(IN1[29]), .S(SEL), .Z(Y[29]) );
  MUX2_X1 U23 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U24 ( .A(IN1[2]), .B(IN1[30]), .S(SEL), .Z(Y[30]) );
  MUX2_X1 U25 ( .A(IN0[31]), .B(IN1[31]), .S(SEL), .Z(Y[31]) );
  MUX2_X1 U26 ( .A(IN0[32]), .B(IN1[32]), .S(SEL), .Z(Y[32]) );
  MUX2_X1 U27 ( .A(IN0[33]), .B(IN1[33]), .S(SEL), .Z(Y[33]) );
  MUX2_X1 U28 ( .A(IN0[34]), .B(IN1[34]), .S(SEL), .Z(Y[34]) );
  MUX2_X1 U29 ( .A(IN0[35]), .B(IN1[35]), .S(SEL), .Z(Y[35]) );
  MUX2_X1 U30 ( .A(IN0[3]), .B(IN0[31]), .S(SEL), .Z(Y[3]) );
  MUX2_X1 U31 ( .A(IN0[4]), .B(IN0[32]), .S(SEL), .Z(Y[4]) );
  MUX2_X1 U32 ( .A(IN0[5]), .B(IN0[33]), .S(SEL), .Z(Y[5]) );
  MUX2_X1 U33 ( .A(IN0[6]), .B(IN0[34]), .S(SEL), .Z(Y[6]) );
  MUX2_X1 U34 ( .A(IN0[7]), .B(IN0[35]), .S(SEL), .Z(Y[7]) );
  MUX2_X1 U35 ( .A(IN0[8]), .B(IN1[8]), .S(SEL), .Z(Y[8]) );
  MUX2_X1 U36 ( .A(IN0[9]), .B(IN1[9]), .S(SEL), .Z(Y[9]) );
endmodule


module MUX_2to1_N36_4 ( IN0, IN1, SEL, Y );
  input [35:0] IN0;
  input [35:0] IN1;
  output [35:0] Y;
  input SEL;
  wire   n8, n9, n10;

  BUF_X2 U1 ( .A(SEL), .Z(n8) );
  BUF_X2 U2 ( .A(SEL), .Z(n10) );
  CLKBUF_X3 U3 ( .A(SEL), .Z(n9) );
  MUX2_X1 U4 ( .A(IN0[21]), .B(IN1[21]), .S(n8), .Z(Y[21]) );
  MUX2_X1 U5 ( .A(IN0[0]), .B(IN1[0]), .S(n9), .Z(Y[0]) );
  MUX2_X1 U6 ( .A(IN0[10]), .B(IN1[10]), .S(n8), .Z(Y[10]) );
  MUX2_X1 U7 ( .A(IN0[11]), .B(IN1[11]), .S(n8), .Z(Y[11]) );
  MUX2_X1 U8 ( .A(IN0[12]), .B(IN1[12]), .S(n8), .Z(Y[12]) );
  MUX2_X1 U9 ( .A(IN0[13]), .B(IN1[13]), .S(n8), .Z(Y[13]) );
  MUX2_X1 U10 ( .A(IN0[14]), .B(IN1[14]), .S(n9), .Z(Y[14]) );
  MUX2_X1 U11 ( .A(IN0[15]), .B(IN1[15]), .S(n8), .Z(Y[15]) );
  MUX2_X1 U12 ( .A(IN0[16]), .B(IN1[16]), .S(n9), .Z(Y[16]) );
  MUX2_X1 U13 ( .A(IN0[17]), .B(IN1[17]), .S(n8), .Z(Y[17]) );
  MUX2_X1 U14 ( .A(IN0[18]), .B(IN1[18]), .S(n8), .Z(Y[18]) );
  MUX2_X1 U15 ( .A(IN0[19]), .B(IN1[19]), .S(n8), .Z(Y[19]) );
  MUX2_X1 U16 ( .A(IN0[1]), .B(IN1[1]), .S(n9), .Z(Y[1]) );
  MUX2_X1 U17 ( .A(IN0[20]), .B(IN1[20]), .S(n10), .Z(Y[20]) );
  MUX2_X1 U18 ( .A(IN0[22]), .B(IN1[22]), .S(n10), .Z(Y[22]) );
  MUX2_X1 U19 ( .A(IN0[23]), .B(IN1[23]), .S(n9), .Z(Y[23]) );
  MUX2_X1 U20 ( .A(IN0[24]), .B(IN1[24]), .S(n10), .Z(Y[24]) );
  MUX2_X1 U21 ( .A(IN0[25]), .B(IN1[25]), .S(n9), .Z(Y[25]) );
  MUX2_X1 U22 ( .A(IN0[26]), .B(IN1[26]), .S(n9), .Z(Y[26]) );
  MUX2_X1 U23 ( .A(IN0[27]), .B(IN1[27]), .S(n9), .Z(Y[27]) );
  MUX2_X1 U24 ( .A(IN0[28]), .B(IN1[28]), .S(n10), .Z(Y[28]) );
  MUX2_X1 U25 ( .A(IN0[29]), .B(IN1[29]), .S(n10), .Z(Y[29]) );
  MUX2_X1 U26 ( .A(IN0[2]), .B(IN1[2]), .S(n10), .Z(Y[2]) );
  MUX2_X1 U27 ( .A(IN0[30]), .B(IN1[30]), .S(n10), .Z(Y[30]) );
  MUX2_X1 U28 ( .A(IN0[31]), .B(IN1[31]), .S(n10), .Z(Y[31]) );
  MUX2_X1 U29 ( .A(IN0[32]), .B(IN1[32]), .S(n9), .Z(Y[32]) );
  MUX2_X1 U30 ( .A(IN0[33]), .B(IN1[33]), .S(n9), .Z(Y[33]) );
  MUX2_X1 U31 ( .A(IN0[34]), .B(IN1[34]), .S(n9), .Z(Y[34]) );
  MUX2_X1 U32 ( .A(IN0[35]), .B(IN1[35]), .S(n10), .Z(Y[35]) );
  MUX2_X1 U33 ( .A(IN0[3]), .B(IN1[3]), .S(n9), .Z(Y[3]) );
  MUX2_X1 U34 ( .A(IN0[4]), .B(IN1[4]), .S(n10), .Z(Y[4]) );
  MUX2_X1 U35 ( .A(IN0[5]), .B(IN1[5]), .S(n9), .Z(Y[5]) );
  MUX2_X1 U36 ( .A(IN0[6]), .B(IN1[6]), .S(n10), .Z(Y[6]) );
  MUX2_X1 U37 ( .A(IN0[7]), .B(IN1[7]), .S(n10), .Z(Y[7]) );
  MUX2_X1 U38 ( .A(IN0[8]), .B(IN1[8]), .S(n10), .Z(Y[8]) );
  MUX2_X1 U39 ( .A(IN0[9]), .B(IN1[9]), .S(n8), .Z(Y[9]) );
endmodule


module MUX_2to1_N36_3 ( IN0, IN1, SEL, Y );
  input [35:0] IN0;
  input [35:0] IN1;
  output [35:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(IN0[10]), .B(IN1[10]), .S(SEL), .Z(Y[10]) );
  MUX2_X1 U3 ( .A(IN0[11]), .B(IN1[11]), .S(SEL), .Z(Y[11]) );
  MUX2_X1 U4 ( .A(IN0[12]), .B(IN1[12]), .S(SEL), .Z(Y[12]) );
  MUX2_X1 U5 ( .A(IN0[13]), .B(IN1[13]), .S(SEL), .Z(Y[13]) );
  MUX2_X1 U6 ( .A(IN0[14]), .B(IN1[14]), .S(SEL), .Z(Y[14]) );
  MUX2_X1 U7 ( .A(IN0[15]), .B(IN1[15]), .S(SEL), .Z(Y[15]) );
  MUX2_X1 U8 ( .A(IN0[16]), .B(IN1[16]), .S(SEL), .Z(Y[16]) );
  MUX2_X1 U9 ( .A(IN0[17]), .B(IN1[17]), .S(SEL), .Z(Y[17]) );
  MUX2_X1 U10 ( .A(IN0[18]), .B(IN1[18]), .S(SEL), .Z(Y[18]) );
  MUX2_X1 U11 ( .A(IN0[19]), .B(IN1[19]), .S(SEL), .Z(Y[19]) );
  MUX2_X1 U12 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U13 ( .A(IN0[20]), .B(IN1[20]), .S(SEL), .Z(Y[20]) );
  MUX2_X1 U14 ( .A(IN0[21]), .B(IN1[21]), .S(SEL), .Z(Y[21]) );
  MUX2_X1 U15 ( .A(IN0[22]), .B(IN1[22]), .S(SEL), .Z(Y[22]) );
  MUX2_X1 U16 ( .A(IN0[23]), .B(IN1[23]), .S(SEL), .Z(Y[23]) );
  MUX2_X1 U17 ( .A(IN0[24]), .B(IN1[24]), .S(SEL), .Z(Y[24]) );
  MUX2_X1 U18 ( .A(IN0[25]), .B(IN1[25]), .S(SEL), .Z(Y[25]) );
  MUX2_X1 U19 ( .A(IN0[26]), .B(IN1[26]), .S(SEL), .Z(Y[26]) );
  MUX2_X1 U20 ( .A(IN0[27]), .B(IN1[27]), .S(SEL), .Z(Y[27]) );
  MUX2_X1 U21 ( .A(IN0[28]), .B(IN1[28]), .S(SEL), .Z(Y[28]) );
  MUX2_X1 U22 ( .A(IN0[29]), .B(IN1[29]), .S(SEL), .Z(Y[29]) );
  MUX2_X1 U23 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U24 ( .A(IN0[30]), .B(IN1[30]), .S(SEL), .Z(Y[30]) );
  MUX2_X1 U25 ( .A(IN0[31]), .B(IN1[31]), .S(SEL), .Z(Y[31]) );
  MUX2_X1 U26 ( .A(IN0[32]), .B(IN1[32]), .S(SEL), .Z(Y[32]) );
  MUX2_X1 U27 ( .A(IN0[33]), .B(IN1[33]), .S(SEL), .Z(Y[33]) );
  MUX2_X1 U28 ( .A(IN0[34]), .B(IN1[34]), .S(SEL), .Z(Y[34]) );
  MUX2_X1 U29 ( .A(IN0[35]), .B(IN1[35]), .S(SEL), .Z(Y[35]) );
  MUX2_X1 U30 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
  MUX2_X1 U31 ( .A(IN0[4]), .B(IN1[4]), .S(SEL), .Z(Y[4]) );
  MUX2_X1 U32 ( .A(IN0[5]), .B(IN1[5]), .S(SEL), .Z(Y[5]) );
  MUX2_X1 U33 ( .A(IN0[6]), .B(IN1[6]), .S(SEL), .Z(Y[6]) );
  MUX2_X1 U34 ( .A(IN0[7]), .B(IN1[7]), .S(SEL), .Z(Y[7]) );
  MUX2_X1 U35 ( .A(IN0[8]), .B(IN1[8]), .S(SEL), .Z(Y[8]) );
  MUX2_X1 U36 ( .A(IN0[9]), .B(IN1[9]), .S(SEL), .Z(Y[9]) );
endmodule


module MUX_2to1_N36_2 ( IN0, IN1, SEL, Y );
  input [35:0] IN0;
  input [35:0] IN1;
  output [35:0] Y;
  input SEL;
  wire   n1, n2, n3, n4, n7, n8, n9;

  AOI22_X1 U1 ( .A1(IN1[9]), .A2(n4), .B1(IN0[9]), .B2(n2), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(Y[9]) );
  CLKBUF_X3 U3 ( .A(SEL), .Z(n8) );
  INV_X1 U4 ( .A(n7), .ZN(n2) );
  INV_X2 U5 ( .A(n2), .ZN(n3) );
  INV_X2 U6 ( .A(n2), .ZN(n4) );
  CLKBUF_X3 U7 ( .A(SEL), .Z(n9) );
  BUF_X1 U8 ( .A(SEL), .Z(n7) );
  MUX2_X1 U9 ( .A(IN0[0]), .B(IN1[0]), .S(n8), .Z(Y[0]) );
  MUX2_X1 U10 ( .A(IN0[10]), .B(IN1[10]), .S(n8), .Z(Y[10]) );
  MUX2_X1 U11 ( .A(IN0[11]), .B(IN1[11]), .S(n8), .Z(Y[11]) );
  MUX2_X1 U12 ( .A(IN0[12]), .B(IN1[12]), .S(n8), .Z(Y[12]) );
  MUX2_X1 U13 ( .A(IN0[13]), .B(IN1[13]), .S(n8), .Z(Y[13]) );
  MUX2_X1 U14 ( .A(IN0[14]), .B(IN1[14]), .S(n8), .Z(Y[14]) );
  MUX2_X1 U15 ( .A(IN0[15]), .B(IN1[15]), .S(n8), .Z(Y[15]) );
  MUX2_X1 U16 ( .A(IN0[16]), .B(IN1[16]), .S(n8), .Z(Y[16]) );
  MUX2_X1 U17 ( .A(IN0[17]), .B(IN1[17]), .S(n8), .Z(Y[17]) );
  MUX2_X1 U18 ( .A(IN0[18]), .B(IN1[18]), .S(n8), .Z(Y[18]) );
  MUX2_X1 U19 ( .A(IN0[19]), .B(IN1[19]), .S(n8), .Z(Y[19]) );
  MUX2_X1 U20 ( .A(IN0[1]), .B(IN1[1]), .S(n9), .Z(Y[1]) );
  MUX2_X1 U21 ( .A(IN0[20]), .B(IN1[20]), .S(n9), .Z(Y[20]) );
  MUX2_X1 U22 ( .A(IN0[21]), .B(IN1[21]), .S(n9), .Z(Y[21]) );
  MUX2_X1 U23 ( .A(IN0[22]), .B(IN1[22]), .S(n9), .Z(Y[22]) );
  MUX2_X1 U24 ( .A(IN0[23]), .B(IN1[23]), .S(n9), .Z(Y[23]) );
  MUX2_X1 U25 ( .A(IN0[24]), .B(IN1[24]), .S(n9), .Z(Y[24]) );
  MUX2_X1 U26 ( .A(IN0[25]), .B(IN1[25]), .S(n9), .Z(Y[25]) );
  MUX2_X1 U27 ( .A(IN0[26]), .B(IN1[26]), .S(n9), .Z(Y[26]) );
  MUX2_X1 U28 ( .A(IN0[27]), .B(IN1[27]), .S(n9), .Z(Y[27]) );
  MUX2_X1 U29 ( .A(IN0[28]), .B(IN1[28]), .S(n9), .Z(Y[28]) );
  MUX2_X1 U30 ( .A(IN0[29]), .B(IN1[29]), .S(n9), .Z(Y[29]) );
  MUX2_X1 U31 ( .A(IN0[2]), .B(IN1[2]), .S(n4), .Z(Y[2]) );
  MUX2_X1 U32 ( .A(IN0[30]), .B(IN1[30]), .S(n4), .Z(Y[30]) );
  MUX2_X1 U33 ( .A(IN0[31]), .B(IN1[31]), .S(n3), .Z(Y[31]) );
  MUX2_X1 U34 ( .A(IN0[32]), .B(IN1[32]), .S(n3), .Z(Y[32]) );
  MUX2_X1 U35 ( .A(IN0[33]), .B(IN1[33]), .S(n3), .Z(Y[33]) );
  MUX2_X1 U36 ( .A(IN0[34]), .B(IN1[34]), .S(n4), .Z(Y[34]) );
  MUX2_X1 U37 ( .A(IN0[35]), .B(IN1[35]), .S(n3), .Z(Y[35]) );
  MUX2_X1 U38 ( .A(IN0[3]), .B(IN1[3]), .S(n4), .Z(Y[3]) );
  MUX2_X1 U39 ( .A(IN0[4]), .B(IN1[4]), .S(n3), .Z(Y[4]) );
  MUX2_X1 U40 ( .A(IN0[5]), .B(IN1[5]), .S(n4), .Z(Y[5]) );
  MUX2_X1 U41 ( .A(IN0[6]), .B(IN1[6]), .S(n3), .Z(Y[6]) );
  MUX2_X1 U42 ( .A(IN0[7]), .B(IN1[7]), .S(n4), .Z(Y[7]) );
  MUX2_X1 U43 ( .A(IN0[8]), .B(IN1[8]), .S(n3), .Z(Y[8]) );
endmodule


module MUX_2to1_N36_1 ( IN0, IN1, SEL, Y );
  input [35:0] IN0;
  input [35:0] IN1;
  output [35:0] Y;
  input SEL;
  wire   n3, n4;

  BUF_X2 U1 ( .A(SEL), .Z(n3) );
  BUF_X2 U2 ( .A(SEL), .Z(n4) );
  MUX2_X1 U3 ( .A(IN0[0]), .B(IN1[0]), .S(n3), .Z(Y[0]) );
  MUX2_X1 U4 ( .A(IN0[10]), .B(IN1[10]), .S(n3), .Z(Y[10]) );
  MUX2_X1 U5 ( .A(IN0[11]), .B(IN1[11]), .S(n3), .Z(Y[11]) );
  MUX2_X1 U6 ( .A(IN0[12]), .B(IN1[12]), .S(n3), .Z(Y[12]) );
  MUX2_X1 U7 ( .A(IN0[13]), .B(IN1[13]), .S(n3), .Z(Y[13]) );
  MUX2_X1 U8 ( .A(IN0[14]), .B(IN1[14]), .S(n3), .Z(Y[14]) );
  MUX2_X1 U9 ( .A(IN0[15]), .B(IN1[15]), .S(n3), .Z(Y[15]) );
  MUX2_X1 U10 ( .A(IN0[16]), .B(IN1[16]), .S(n3), .Z(Y[16]) );
  MUX2_X1 U11 ( .A(IN0[17]), .B(IN1[17]), .S(n3), .Z(Y[17]) );
  MUX2_X1 U12 ( .A(IN0[18]), .B(IN1[18]), .S(n3), .Z(Y[18]) );
  MUX2_X1 U13 ( .A(IN0[19]), .B(IN1[19]), .S(n3), .Z(Y[19]) );
  MUX2_X1 U14 ( .A(IN0[1]), .B(IN1[1]), .S(n3), .Z(Y[1]) );
  MUX2_X1 U15 ( .A(IN0[20]), .B(IN1[20]), .S(SEL), .Z(Y[20]) );
  MUX2_X1 U16 ( .A(IN0[21]), .B(IN1[21]), .S(n4), .Z(Y[21]) );
  MUX2_X1 U17 ( .A(IN0[22]), .B(IN1[22]), .S(n4), .Z(Y[22]) );
  MUX2_X1 U18 ( .A(IN0[23]), .B(IN1[23]), .S(SEL), .Z(Y[23]) );
  MUX2_X1 U19 ( .A(IN0[24]), .B(IN1[24]), .S(SEL), .Z(Y[24]) );
  MUX2_X1 U20 ( .A(IN0[25]), .B(IN1[25]), .S(SEL), .Z(Y[25]) );
  MUX2_X1 U21 ( .A(IN0[26]), .B(IN1[26]), .S(n3), .Z(Y[26]) );
  MUX2_X1 U22 ( .A(IN0[27]), .B(IN1[27]), .S(SEL), .Z(Y[27]) );
  MUX2_X1 U23 ( .A(IN0[28]), .B(IN1[28]), .S(SEL), .Z(Y[28]) );
  MUX2_X1 U24 ( .A(IN0[29]), .B(IN1[29]), .S(SEL), .Z(Y[29]) );
  MUX2_X1 U25 ( .A(IN0[2]), .B(IN1[2]), .S(n4), .Z(Y[2]) );
  MUX2_X1 U26 ( .A(IN0[30]), .B(IN1[30]), .S(n4), .Z(Y[30]) );
  MUX2_X1 U27 ( .A(IN0[31]), .B(IN1[31]), .S(n4), .Z(Y[31]) );
  MUX2_X1 U28 ( .A(IN0[32]), .B(IN1[32]), .S(n4), .Z(Y[32]) );
  MUX2_X1 U29 ( .A(IN0[33]), .B(IN1[33]), .S(n4), .Z(Y[33]) );
  MUX2_X1 U30 ( .A(IN0[34]), .B(IN1[34]), .S(n4), .Z(Y[34]) );
  MUX2_X1 U31 ( .A(IN0[35]), .B(IN1[35]), .S(n4), .Z(Y[35]) );
  MUX2_X1 U32 ( .A(IN0[3]), .B(IN1[3]), .S(n4), .Z(Y[3]) );
  MUX2_X1 U33 ( .A(IN0[4]), .B(IN1[4]), .S(n4), .Z(Y[4]) );
  MUX2_X1 U34 ( .A(IN0[5]), .B(IN1[5]), .S(n4), .Z(Y[5]) );
  MUX2_X1 U35 ( .A(IN0[6]), .B(IN1[6]), .S(n4), .Z(Y[6]) );
  MUX2_X1 U36 ( .A(IN0[7]), .B(IN1[7]), .S(SEL), .Z(Y[7]) );
  MUX2_X1 U37 ( .A(IN0[8]), .B(IN1[8]), .S(SEL), .Z(Y[8]) );
  MUX2_X1 U38 ( .A(IN0[9]), .B(IN1[9]), .S(SEL), .Z(Y[9]) );
endmodule


module MUX_8to1_N36 ( IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, SEL, Y );
  input [35:0] IN0;
  input [35:0] IN1;
  input [35:0] IN2;
  input [35:0] IN3;
  input [35:0] IN4;
  input [35:0] IN5;
  input [35:0] IN6;
  input [35:0] IN7;
  input [2:0] SEL;
  output [35:0] Y;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164;

  AOI22_X1 U1 ( .A1(IN5[10]), .A2(n6), .B1(IN4[10]), .B2(n5), .ZN(n1) );
  AOI22_X1 U2 ( .A1(IN7[10]), .A2(n7), .B1(IN6[10]), .B2(n4), .ZN(n2) );
  NAND4_X1 U3 ( .A1(n20), .A2(n19), .A3(n1), .A4(n2), .ZN(Y[10]) );
  BUF_X2 U4 ( .A(n155), .Z(n3) );
  BUF_X2 U5 ( .A(n160), .Z(n4) );
  BUF_X2 U6 ( .A(n158), .Z(n5) );
  BUF_X2 U7 ( .A(n157), .Z(n6) );
  BUF_X2 U8 ( .A(n159), .Z(n7) );
  BUF_X2 U9 ( .A(n153), .Z(n8) );
  BUF_X2 U10 ( .A(n156), .Z(n9) );
  BUF_X2 U11 ( .A(n154), .Z(n10) );
  NOR3_X1 U12 ( .A1(SEL[2]), .A2(SEL[0]), .A3(SEL[1]), .ZN(n154) );
  INV_X1 U13 ( .A(SEL[0]), .ZN(n11) );
  NOR3_X1 U14 ( .A1(SEL[2]), .A2(SEL[1]), .A3(n11), .ZN(n153) );
  AOI22_X1 U15 ( .A1(n10), .A2(IN0[0]), .B1(n8), .B2(IN1[0]), .ZN(n18) );
  INV_X1 U16 ( .A(SEL[1]), .ZN(n12) );
  NOR3_X1 U17 ( .A1(SEL[2]), .A2(SEL[0]), .A3(n12), .ZN(n156) );
  NAND2_X1 U18 ( .A1(SEL[0]), .A2(SEL[1]), .ZN(n13) );
  NOR2_X1 U19 ( .A1(SEL[2]), .A2(n13), .ZN(n155) );
  AOI22_X1 U20 ( .A1(n9), .A2(IN2[0]), .B1(n155), .B2(IN3[0]), .ZN(n17) );
  INV_X1 U21 ( .A(SEL[2]), .ZN(n14) );
  NOR3_X1 U22 ( .A1(SEL[0]), .A2(SEL[1]), .A3(n14), .ZN(n158) );
  NOR3_X1 U23 ( .A1(SEL[1]), .A2(n11), .A3(n14), .ZN(n157) );
  AOI22_X1 U24 ( .A1(n5), .A2(IN4[0]), .B1(n6), .B2(IN5[0]), .ZN(n16) );
  NOR3_X1 U25 ( .A1(SEL[0]), .A2(n14), .A3(n12), .ZN(n160) );
  NOR2_X1 U26 ( .A1(n14), .A2(n13), .ZN(n159) );
  AOI22_X1 U27 ( .A1(n4), .A2(IN6[0]), .B1(n159), .B2(IN7[0]), .ZN(n15) );
  NAND4_X1 U28 ( .A1(n18), .A2(n17), .A3(n16), .A4(n15), .ZN(Y[0]) );
  AOI22_X1 U29 ( .A1(n10), .A2(IN0[10]), .B1(n8), .B2(IN1[10]), .ZN(n20) );
  AOI22_X1 U30 ( .A1(n9), .A2(IN2[10]), .B1(n3), .B2(IN3[10]), .ZN(n19) );
  AOI22_X1 U31 ( .A1(n10), .A2(IN0[11]), .B1(n8), .B2(IN1[11]), .ZN(n24) );
  AOI22_X1 U32 ( .A1(n9), .A2(IN2[11]), .B1(n155), .B2(IN3[11]), .ZN(n23) );
  AOI22_X1 U33 ( .A1(n5), .A2(IN4[11]), .B1(n6), .B2(IN5[11]), .ZN(n22) );
  AOI22_X1 U34 ( .A1(n4), .A2(IN6[11]), .B1(n159), .B2(IN7[11]), .ZN(n21) );
  NAND4_X1 U35 ( .A1(n24), .A2(n23), .A3(n22), .A4(n21), .ZN(Y[11]) );
  AOI22_X1 U36 ( .A1(n10), .A2(IN0[12]), .B1(n8), .B2(IN1[12]), .ZN(n28) );
  AOI22_X1 U37 ( .A1(n9), .A2(IN2[12]), .B1(n3), .B2(IN3[12]), .ZN(n27) );
  AOI22_X1 U38 ( .A1(n5), .A2(IN4[12]), .B1(n6), .B2(IN5[12]), .ZN(n26) );
  AOI22_X1 U39 ( .A1(n4), .A2(IN6[12]), .B1(n7), .B2(IN7[12]), .ZN(n25) );
  NAND4_X1 U40 ( .A1(n28), .A2(n27), .A3(n26), .A4(n25), .ZN(Y[12]) );
  AOI22_X1 U41 ( .A1(n10), .A2(IN0[13]), .B1(n153), .B2(IN1[13]), .ZN(n32) );
  AOI22_X1 U42 ( .A1(n9), .A2(IN2[13]), .B1(n155), .B2(IN3[13]), .ZN(n31) );
  AOI22_X1 U43 ( .A1(n5), .A2(IN4[13]), .B1(n157), .B2(IN5[13]), .ZN(n30) );
  AOI22_X1 U44 ( .A1(n4), .A2(IN6[13]), .B1(n159), .B2(IN7[13]), .ZN(n29) );
  NAND4_X1 U45 ( .A1(n32), .A2(n31), .A3(n30), .A4(n29), .ZN(Y[13]) );
  AOI22_X1 U46 ( .A1(n10), .A2(IN0[14]), .B1(n8), .B2(IN1[14]), .ZN(n36) );
  AOI22_X1 U47 ( .A1(n9), .A2(IN2[14]), .B1(n3), .B2(IN3[14]), .ZN(n35) );
  AOI22_X1 U48 ( .A1(n5), .A2(IN4[14]), .B1(n6), .B2(IN5[14]), .ZN(n34) );
  AOI22_X1 U49 ( .A1(n4), .A2(IN6[14]), .B1(n7), .B2(IN7[14]), .ZN(n33) );
  NAND4_X1 U50 ( .A1(n36), .A2(n35), .A3(n34), .A4(n33), .ZN(Y[14]) );
  AOI22_X1 U51 ( .A1(n10), .A2(IN0[15]), .B1(n153), .B2(IN1[15]), .ZN(n40) );
  AOI22_X1 U52 ( .A1(n9), .A2(IN2[15]), .B1(n155), .B2(IN3[15]), .ZN(n39) );
  AOI22_X1 U53 ( .A1(n5), .A2(IN4[15]), .B1(n157), .B2(IN5[15]), .ZN(n38) );
  AOI22_X1 U54 ( .A1(n4), .A2(IN6[15]), .B1(n159), .B2(IN7[15]), .ZN(n37) );
  NAND4_X1 U55 ( .A1(n40), .A2(n39), .A3(n38), .A4(n37), .ZN(Y[15]) );
  AOI22_X1 U56 ( .A1(n10), .A2(IN0[16]), .B1(n8), .B2(IN1[16]), .ZN(n44) );
  AOI22_X1 U57 ( .A1(n9), .A2(IN2[16]), .B1(n3), .B2(IN3[16]), .ZN(n43) );
  AOI22_X1 U58 ( .A1(n5), .A2(IN4[16]), .B1(n6), .B2(IN5[16]), .ZN(n42) );
  AOI22_X1 U59 ( .A1(n4), .A2(IN6[16]), .B1(n7), .B2(IN7[16]), .ZN(n41) );
  NAND4_X1 U60 ( .A1(n44), .A2(n43), .A3(n42), .A4(n41), .ZN(Y[16]) );
  AOI22_X1 U61 ( .A1(n10), .A2(IN0[17]), .B1(n153), .B2(IN1[17]), .ZN(n48) );
  AOI22_X1 U62 ( .A1(n9), .A2(IN2[17]), .B1(n155), .B2(IN3[17]), .ZN(n47) );
  AOI22_X1 U63 ( .A1(n5), .A2(IN4[17]), .B1(n157), .B2(IN5[17]), .ZN(n46) );
  AOI22_X1 U64 ( .A1(n4), .A2(IN6[17]), .B1(n159), .B2(IN7[17]), .ZN(n45) );
  NAND4_X1 U65 ( .A1(n45), .A2(n47), .A3(n46), .A4(n48), .ZN(Y[17]) );
  AOI22_X1 U66 ( .A1(n10), .A2(IN0[18]), .B1(n8), .B2(IN1[18]), .ZN(n52) );
  AOI22_X1 U67 ( .A1(n9), .A2(IN2[18]), .B1(n3), .B2(IN3[18]), .ZN(n51) );
  AOI22_X1 U68 ( .A1(n5), .A2(IN4[18]), .B1(n6), .B2(IN5[18]), .ZN(n50) );
  AOI22_X1 U69 ( .A1(n4), .A2(IN6[18]), .B1(n7), .B2(IN7[18]), .ZN(n49) );
  NAND4_X1 U70 ( .A1(n52), .A2(n51), .A3(n50), .A4(n49), .ZN(Y[18]) );
  AOI22_X1 U71 ( .A1(n10), .A2(IN0[19]), .B1(n153), .B2(IN1[19]), .ZN(n56) );
  AOI22_X1 U72 ( .A1(n9), .A2(IN2[19]), .B1(n155), .B2(IN3[19]), .ZN(n55) );
  AOI22_X1 U73 ( .A1(n5), .A2(IN4[19]), .B1(n157), .B2(IN5[19]), .ZN(n54) );
  AOI22_X1 U74 ( .A1(n4), .A2(IN6[19]), .B1(n159), .B2(IN7[19]), .ZN(n53) );
  NAND4_X1 U75 ( .A1(n56), .A2(n55), .A3(n54), .A4(n53), .ZN(Y[19]) );
  AOI22_X1 U76 ( .A1(n10), .A2(IN0[1]), .B1(n8), .B2(IN1[1]), .ZN(n60) );
  AOI22_X1 U77 ( .A1(n9), .A2(IN2[1]), .B1(n3), .B2(IN3[1]), .ZN(n59) );
  AOI22_X1 U78 ( .A1(n5), .A2(IN4[1]), .B1(n6), .B2(IN5[1]), .ZN(n58) );
  AOI22_X1 U79 ( .A1(n4), .A2(IN6[1]), .B1(n7), .B2(IN7[1]), .ZN(n57) );
  NAND4_X1 U80 ( .A1(n60), .A2(n59), .A3(n58), .A4(n57), .ZN(Y[1]) );
  AOI22_X1 U81 ( .A1(n10), .A2(IN0[20]), .B1(n8), .B2(IN1[20]), .ZN(n64) );
  AOI22_X1 U82 ( .A1(n9), .A2(IN2[20]), .B1(n3), .B2(IN3[20]), .ZN(n63) );
  AOI22_X1 U83 ( .A1(n5), .A2(IN4[20]), .B1(n6), .B2(IN5[20]), .ZN(n62) );
  AOI22_X1 U84 ( .A1(n4), .A2(IN6[20]), .B1(n7), .B2(IN7[20]), .ZN(n61) );
  NAND4_X1 U85 ( .A1(n64), .A2(n63), .A3(n62), .A4(n61), .ZN(Y[20]) );
  AOI22_X1 U86 ( .A1(n10), .A2(IN0[21]), .B1(n8), .B2(IN1[21]), .ZN(n68) );
  AOI22_X1 U87 ( .A1(n9), .A2(IN2[21]), .B1(n3), .B2(IN3[21]), .ZN(n67) );
  AOI22_X1 U88 ( .A1(n5), .A2(IN4[21]), .B1(n6), .B2(IN5[21]), .ZN(n66) );
  AOI22_X1 U89 ( .A1(n4), .A2(IN6[21]), .B1(n7), .B2(IN7[21]), .ZN(n65) );
  NAND4_X1 U90 ( .A1(n68), .A2(n67), .A3(n66), .A4(n65), .ZN(Y[21]) );
  AOI22_X1 U91 ( .A1(n10), .A2(IN0[22]), .B1(n8), .B2(IN1[22]), .ZN(n72) );
  AOI22_X1 U92 ( .A1(n9), .A2(IN2[22]), .B1(n3), .B2(IN3[22]), .ZN(n71) );
  AOI22_X1 U93 ( .A1(n5), .A2(IN4[22]), .B1(n6), .B2(IN5[22]), .ZN(n70) );
  AOI22_X1 U94 ( .A1(n4), .A2(IN6[22]), .B1(n7), .B2(IN7[22]), .ZN(n69) );
  NAND4_X1 U95 ( .A1(n72), .A2(n71), .A3(n70), .A4(n69), .ZN(Y[22]) );
  AOI22_X1 U96 ( .A1(n10), .A2(IN0[23]), .B1(n8), .B2(IN1[23]), .ZN(n76) );
  AOI22_X1 U97 ( .A1(n9), .A2(IN2[23]), .B1(n3), .B2(IN3[23]), .ZN(n75) );
  AOI22_X1 U98 ( .A1(n5), .A2(IN4[23]), .B1(n6), .B2(IN5[23]), .ZN(n74) );
  AOI22_X1 U99 ( .A1(n4), .A2(IN6[23]), .B1(n7), .B2(IN7[23]), .ZN(n73) );
  NAND4_X1 U100 ( .A1(n76), .A2(n75), .A3(n74), .A4(n73), .ZN(Y[23]) );
  AOI22_X1 U101 ( .A1(n10), .A2(IN0[24]), .B1(n8), .B2(IN1[24]), .ZN(n80) );
  AOI22_X1 U102 ( .A1(n9), .A2(IN2[24]), .B1(n3), .B2(IN3[24]), .ZN(n79) );
  AOI22_X1 U103 ( .A1(n5), .A2(IN4[24]), .B1(n6), .B2(IN5[24]), .ZN(n78) );
  AOI22_X1 U104 ( .A1(n4), .A2(IN6[24]), .B1(n7), .B2(IN7[24]), .ZN(n77) );
  NAND4_X1 U105 ( .A1(n80), .A2(n79), .A3(n78), .A4(n77), .ZN(Y[24]) );
  AOI22_X1 U106 ( .A1(n10), .A2(IN0[25]), .B1(n8), .B2(IN1[25]), .ZN(n84) );
  AOI22_X1 U107 ( .A1(n9), .A2(IN2[25]), .B1(n155), .B2(IN3[25]), .ZN(n83) );
  AOI22_X1 U108 ( .A1(n5), .A2(IN4[25]), .B1(n6), .B2(IN5[25]), .ZN(n82) );
  AOI22_X1 U109 ( .A1(n4), .A2(IN6[25]), .B1(n159), .B2(IN7[25]), .ZN(n81) );
  NAND4_X1 U110 ( .A1(n84), .A2(n83), .A3(n82), .A4(n81), .ZN(Y[25]) );
  AOI22_X1 U111 ( .A1(n10), .A2(IN0[26]), .B1(n8), .B2(IN1[26]), .ZN(n88) );
  AOI22_X1 U112 ( .A1(n9), .A2(IN2[26]), .B1(n3), .B2(IN3[26]), .ZN(n87) );
  AOI22_X1 U113 ( .A1(n5), .A2(IN4[26]), .B1(n6), .B2(IN5[26]), .ZN(n86) );
  AOI22_X1 U114 ( .A1(n4), .A2(IN6[26]), .B1(n7), .B2(IN7[26]), .ZN(n85) );
  NAND4_X1 U115 ( .A1(n88), .A2(n87), .A3(n86), .A4(n85), .ZN(Y[26]) );
  AOI22_X1 U116 ( .A1(n10), .A2(IN0[27]), .B1(n8), .B2(IN1[27]), .ZN(n92) );
  AOI22_X1 U117 ( .A1(n9), .A2(IN2[27]), .B1(n155), .B2(IN3[27]), .ZN(n91) );
  AOI22_X1 U118 ( .A1(n5), .A2(IN4[27]), .B1(n6), .B2(IN5[27]), .ZN(n90) );
  AOI22_X1 U119 ( .A1(n4), .A2(IN6[27]), .B1(n159), .B2(IN7[27]), .ZN(n89) );
  NAND4_X1 U120 ( .A1(n92), .A2(n91), .A3(n90), .A4(n89), .ZN(Y[27]) );
  AOI22_X1 U121 ( .A1(n10), .A2(IN0[28]), .B1(n8), .B2(IN1[28]), .ZN(n96) );
  AOI22_X1 U122 ( .A1(n9), .A2(IN2[28]), .B1(n3), .B2(IN3[28]), .ZN(n95) );
  AOI22_X1 U123 ( .A1(n5), .A2(IN4[28]), .B1(n6), .B2(IN5[28]), .ZN(n94) );
  AOI22_X1 U124 ( .A1(n4), .A2(IN6[28]), .B1(n7), .B2(IN7[28]), .ZN(n93) );
  NAND4_X1 U125 ( .A1(n96), .A2(n95), .A3(n94), .A4(n93), .ZN(Y[28]) );
  AOI22_X1 U126 ( .A1(n10), .A2(IN0[29]), .B1(n153), .B2(IN1[29]), .ZN(n100)
         );
  AOI22_X1 U127 ( .A1(n9), .A2(IN2[29]), .B1(n155), .B2(IN3[29]), .ZN(n99) );
  AOI22_X1 U128 ( .A1(n5), .A2(IN4[29]), .B1(n157), .B2(IN5[29]), .ZN(n98) );
  AOI22_X1 U129 ( .A1(n4), .A2(IN6[29]), .B1(n159), .B2(IN7[29]), .ZN(n97) );
  NAND4_X1 U130 ( .A1(n100), .A2(n99), .A3(n98), .A4(n97), .ZN(Y[29]) );
  AOI22_X1 U131 ( .A1(n10), .A2(IN0[2]), .B1(n8), .B2(IN1[2]), .ZN(n104) );
  AOI22_X1 U132 ( .A1(n9), .A2(IN2[2]), .B1(n3), .B2(IN3[2]), .ZN(n103) );
  AOI22_X1 U133 ( .A1(n5), .A2(IN4[2]), .B1(n6), .B2(IN5[2]), .ZN(n102) );
  AOI22_X1 U134 ( .A1(n4), .A2(IN6[2]), .B1(n7), .B2(IN7[2]), .ZN(n101) );
  NAND4_X1 U135 ( .A1(n104), .A2(n103), .A3(n102), .A4(n101), .ZN(Y[2]) );
  AOI22_X1 U136 ( .A1(n154), .A2(IN0[30]), .B1(n8), .B2(IN1[30]), .ZN(n108) );
  AOI22_X1 U137 ( .A1(n156), .A2(IN2[30]), .B1(n3), .B2(IN3[30]), .ZN(n107) );
  AOI22_X1 U138 ( .A1(n158), .A2(IN4[30]), .B1(n6), .B2(IN5[30]), .ZN(n106) );
  AOI22_X1 U139 ( .A1(n160), .A2(IN6[30]), .B1(n7), .B2(IN7[30]), .ZN(n105) );
  NAND4_X1 U140 ( .A1(n108), .A2(n107), .A3(n106), .A4(n105), .ZN(Y[30]) );
  AOI22_X1 U141 ( .A1(n154), .A2(IN0[31]), .B1(n8), .B2(IN1[31]), .ZN(n112) );
  AOI22_X1 U142 ( .A1(n156), .A2(IN2[31]), .B1(n3), .B2(IN3[31]), .ZN(n111) );
  AOI22_X1 U143 ( .A1(n158), .A2(IN4[31]), .B1(n6), .B2(IN5[31]), .ZN(n110) );
  AOI22_X1 U144 ( .A1(n160), .A2(IN6[31]), .B1(n7), .B2(IN7[31]), .ZN(n109) );
  NAND4_X1 U145 ( .A1(n112), .A2(n111), .A3(n110), .A4(n109), .ZN(Y[31]) );
  AOI22_X1 U146 ( .A1(n10), .A2(IN0[32]), .B1(n8), .B2(IN1[32]), .ZN(n116) );
  AOI22_X1 U147 ( .A1(n9), .A2(IN2[32]), .B1(n3), .B2(IN3[32]), .ZN(n115) );
  AOI22_X1 U148 ( .A1(n5), .A2(IN4[32]), .B1(n6), .B2(IN5[32]), .ZN(n114) );
  AOI22_X1 U149 ( .A1(n4), .A2(IN6[32]), .B1(n7), .B2(IN7[32]), .ZN(n113) );
  NAND4_X1 U150 ( .A1(n116), .A2(n115), .A3(n114), .A4(n113), .ZN(Y[32]) );
  AOI22_X1 U151 ( .A1(n154), .A2(IN0[33]), .B1(n8), .B2(IN1[33]), .ZN(n120) );
  AOI22_X1 U152 ( .A1(n156), .A2(IN2[33]), .B1(n3), .B2(IN3[33]), .ZN(n119) );
  AOI22_X1 U153 ( .A1(n158), .A2(IN4[33]), .B1(n6), .B2(IN5[33]), .ZN(n118) );
  AOI22_X1 U154 ( .A1(n160), .A2(IN6[33]), .B1(n7), .B2(IN7[33]), .ZN(n117) );
  NAND4_X1 U155 ( .A1(n120), .A2(n119), .A3(n118), .A4(n117), .ZN(Y[33]) );
  AOI22_X1 U156 ( .A1(n10), .A2(IN0[34]), .B1(n8), .B2(IN1[34]), .ZN(n124) );
  AOI22_X1 U157 ( .A1(n9), .A2(IN2[34]), .B1(n3), .B2(IN3[34]), .ZN(n123) );
  AOI22_X1 U158 ( .A1(n5), .A2(IN4[34]), .B1(n6), .B2(IN5[34]), .ZN(n122) );
  AOI22_X1 U159 ( .A1(n4), .A2(IN6[34]), .B1(n7), .B2(IN7[34]), .ZN(n121) );
  NAND4_X1 U160 ( .A1(n124), .A2(n123), .A3(n122), .A4(n121), .ZN(Y[34]) );
  AOI22_X1 U161 ( .A1(n10), .A2(IN0[35]), .B1(n8), .B2(IN1[35]), .ZN(n128) );
  AOI22_X1 U162 ( .A1(n9), .A2(IN2[35]), .B1(n3), .B2(IN3[35]), .ZN(n127) );
  AOI22_X1 U163 ( .A1(n5), .A2(IN4[35]), .B1(n6), .B2(IN5[35]), .ZN(n126) );
  AOI22_X1 U164 ( .A1(n4), .A2(IN6[35]), .B1(n7), .B2(IN7[35]), .ZN(n125) );
  NAND4_X1 U165 ( .A1(n128), .A2(n127), .A3(n126), .A4(n125), .ZN(Y[35]) );
  AOI22_X1 U166 ( .A1(n154), .A2(IN0[3]), .B1(n8), .B2(IN1[3]), .ZN(n132) );
  AOI22_X1 U167 ( .A1(n156), .A2(IN2[3]), .B1(n3), .B2(IN3[3]), .ZN(n131) );
  AOI22_X1 U168 ( .A1(n158), .A2(IN4[3]), .B1(n6), .B2(IN5[3]), .ZN(n130) );
  AOI22_X1 U169 ( .A1(n160), .A2(IN6[3]), .B1(n7), .B2(IN7[3]), .ZN(n129) );
  NAND4_X1 U170 ( .A1(n132), .A2(n131), .A3(n130), .A4(n129), .ZN(Y[3]) );
  AOI22_X1 U171 ( .A1(n10), .A2(IN0[4]), .B1(n8), .B2(IN1[4]), .ZN(n136) );
  AOI22_X1 U172 ( .A1(n9), .A2(IN2[4]), .B1(n3), .B2(IN3[4]), .ZN(n135) );
  AOI22_X1 U173 ( .A1(n5), .A2(IN4[4]), .B1(n6), .B2(IN5[4]), .ZN(n134) );
  AOI22_X1 U174 ( .A1(n4), .A2(IN6[4]), .B1(n7), .B2(IN7[4]), .ZN(n133) );
  NAND4_X1 U175 ( .A1(n136), .A2(n135), .A3(n134), .A4(n133), .ZN(Y[4]) );
  AOI22_X1 U176 ( .A1(n154), .A2(IN0[5]), .B1(n8), .B2(IN1[5]), .ZN(n140) );
  AOI22_X1 U177 ( .A1(n156), .A2(IN2[5]), .B1(n3), .B2(IN3[5]), .ZN(n139) );
  AOI22_X1 U178 ( .A1(n158), .A2(IN4[5]), .B1(n6), .B2(IN5[5]), .ZN(n138) );
  AOI22_X1 U179 ( .A1(n160), .A2(IN6[5]), .B1(n7), .B2(IN7[5]), .ZN(n137) );
  NAND4_X1 U180 ( .A1(n140), .A2(n139), .A3(n138), .A4(n137), .ZN(Y[5]) );
  AOI22_X1 U181 ( .A1(n10), .A2(IN0[6]), .B1(n8), .B2(IN1[6]), .ZN(n144) );
  AOI22_X1 U182 ( .A1(n9), .A2(IN2[6]), .B1(n3), .B2(IN3[6]), .ZN(n143) );
  AOI22_X1 U183 ( .A1(n5), .A2(IN4[6]), .B1(n6), .B2(IN5[6]), .ZN(n142) );
  AOI22_X1 U184 ( .A1(n4), .A2(IN6[6]), .B1(n7), .B2(IN7[6]), .ZN(n141) );
  NAND4_X1 U185 ( .A1(n144), .A2(n143), .A3(n142), .A4(n141), .ZN(Y[6]) );
  AOI22_X1 U186 ( .A1(n10), .A2(IN0[7]), .B1(n8), .B2(IN1[7]), .ZN(n148) );
  AOI22_X1 U187 ( .A1(n9), .A2(IN2[7]), .B1(n3), .B2(IN3[7]), .ZN(n147) );
  AOI22_X1 U188 ( .A1(n5), .A2(IN4[7]), .B1(n6), .B2(IN5[7]), .ZN(n146) );
  AOI22_X1 U189 ( .A1(n4), .A2(IN6[7]), .B1(n7), .B2(IN7[7]), .ZN(n145) );
  NAND4_X1 U190 ( .A1(n148), .A2(n147), .A3(n146), .A4(n145), .ZN(Y[7]) );
  AOI22_X1 U191 ( .A1(n10), .A2(IN0[8]), .B1(n8), .B2(IN1[8]), .ZN(n152) );
  AOI22_X1 U192 ( .A1(n9), .A2(IN2[8]), .B1(n3), .B2(IN3[8]), .ZN(n151) );
  AOI22_X1 U193 ( .A1(n5), .A2(IN4[8]), .B1(n6), .B2(IN5[8]), .ZN(n150) );
  AOI22_X1 U194 ( .A1(n4), .A2(IN6[8]), .B1(n7), .B2(IN7[8]), .ZN(n149) );
  NAND4_X1 U195 ( .A1(n152), .A2(n151), .A3(n150), .A4(n149), .ZN(Y[8]) );
  AOI22_X1 U196 ( .A1(n10), .A2(IN0[9]), .B1(n8), .B2(IN1[9]), .ZN(n164) );
  AOI22_X1 U197 ( .A1(n9), .A2(IN2[9]), .B1(n3), .B2(IN3[9]), .ZN(n163) );
  AOI22_X1 U198 ( .A1(n5), .A2(IN4[9]), .B1(n6), .B2(IN5[9]), .ZN(n162) );
  AOI22_X1 U199 ( .A1(n4), .A2(IN6[9]), .B1(n7), .B2(IN7[9]), .ZN(n161) );
  NAND4_X1 U200 ( .A1(n164), .A2(n163), .A3(n162), .A4(n161), .ZN(Y[9]) );
endmodule


module MUX_8to1_N32_1 ( IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, SEL, Y );
  input [31:0] IN0;
  input [31:0] IN1;
  input [31:0] IN2;
  input [31:0] IN3;
  input [31:0] IN4;
  input [31:0] IN5;
  input [31:0] IN6;
  input [31:0] IN7;
  input [2:0] SEL;
  output [31:0] Y;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98;

  OR2_X1 U1 ( .A1(n36), .A2(n98), .ZN(n4) );
  OR2_X1 U2 ( .A1(n36), .A2(n91), .ZN(n5) );
  OAI211_X1 U3 ( .C1(n26), .C2(n98), .A(n23), .B(n22), .ZN(Y[13]) );
  INV_X2 U4 ( .A(n91), .ZN(n94) );
  INV_X1 U5 ( .A(n87), .ZN(n98) );
  INV_X2 U6 ( .A(n7), .ZN(n1) );
  OR2_X1 U7 ( .A1(n21), .A2(n98), .ZN(n3) );
  BUF_X2 U8 ( .A(n92), .Z(n2) );
  NAND3_X1 U9 ( .A1(n19), .A2(n20), .A3(n3), .ZN(Y[12]) );
  NAND3_X1 U10 ( .A1(n33), .A2(n32), .A3(n4), .ZN(Y[17]) );
  NAND3_X1 U11 ( .A1(n34), .A2(n35), .A3(n5), .ZN(Y[18]) );
  BUF_X1 U12 ( .A(IN0[3]), .Z(n6) );
  OR2_X1 U13 ( .A1(n11), .A2(n9), .ZN(n7) );
  NOR2_X2 U14 ( .A1(n10), .A2(n11), .ZN(n87) );
  BUF_X1 U15 ( .A(n93), .Z(n8) );
  INV_X1 U16 ( .A(SEL[0]), .ZN(n11) );
  XOR2_X1 U17 ( .A(SEL[1]), .B(SEL[2]), .Z(n9) );
  INV_X1 U18 ( .A(IN7[0]), .ZN(n68) );
  INV_X1 U19 ( .A(SEL[1]), .ZN(n12) );
  NOR2_X1 U20 ( .A1(SEL[0]), .A2(n12), .ZN(n93) );
  NOR3_X1 U21 ( .A1(SEL[1]), .A2(SEL[2]), .A3(SEL[0]), .ZN(n92) );
  AOI22_X1 U22 ( .A1(n8), .A2(IN6[0]), .B1(n2), .B2(IN0[0]), .ZN(n14) );
  INV_X1 U23 ( .A(n9), .ZN(n10) );
  NAND3_X1 U24 ( .A1(n12), .A2(n11), .A3(SEL[2]), .ZN(n91) );
  AOI22_X1 U25 ( .A1(n87), .A2(IN5[0]), .B1(n94), .B2(IN4[0]), .ZN(n13) );
  OAI211_X1 U26 ( .C1(n7), .C2(n68), .A(n14), .B(n13), .ZN(Y[0]) );
  INV_X1 U27 ( .A(IN7[10]), .ZN(n21) );
  AOI22_X1 U28 ( .A1(n8), .A2(IN6[10]), .B1(n2), .B2(IN0[10]), .ZN(n16) );
  AOI22_X1 U29 ( .A1(n87), .A2(IN5[10]), .B1(n94), .B2(IN4[10]), .ZN(n15) );
  OAI211_X1 U30 ( .C1(n7), .C2(n21), .A(n16), .B(n15), .ZN(Y[10]) );
  INV_X1 U31 ( .A(IN0[10]), .ZN(n26) );
  AOI22_X1 U32 ( .A1(n8), .A2(IN7[10]), .B1(n2), .B2(IN0[11]), .ZN(n18) );
  AOI22_X1 U33 ( .A1(n87), .A2(IN6[10]), .B1(IN5[10]), .B2(n94), .ZN(n17) );
  OAI211_X1 U34 ( .C1(n7), .C2(n26), .A(n17), .B(n18), .ZN(Y[11]) );
  AOI22_X1 U35 ( .A1(n8), .A2(IN0[10]), .B1(n2), .B2(IN0[12]), .ZN(n20) );
  AOI22_X1 U36 ( .A1(n1), .A2(IN0[11]), .B1(n94), .B2(IN6[10]), .ZN(n19) );
  AOI22_X1 U37 ( .A1(n8), .A2(IN0[11]), .B1(n2), .B2(IN0[13]), .ZN(n23) );
  AOI22_X1 U38 ( .A1(n1), .A2(IN0[12]), .B1(n94), .B2(IN7[10]), .ZN(n22) );
  AOI22_X1 U39 ( .A1(n8), .A2(IN0[12]), .B1(n2), .B2(IN0[14]), .ZN(n25) );
  AOI22_X1 U40 ( .A1(n87), .A2(IN0[11]), .B1(n1), .B2(IN0[13]), .ZN(n24) );
  OAI211_X1 U41 ( .C1(n91), .C2(n26), .A(n25), .B(n24), .ZN(Y[14]) );
  INV_X1 U42 ( .A(IN0[12]), .ZN(n31) );
  AOI22_X1 U43 ( .A1(n8), .A2(IN0[13]), .B1(n2), .B2(IN0[15]), .ZN(n28) );
  AOI22_X1 U44 ( .A1(n1), .A2(IN0[14]), .B1(n94), .B2(IN0[11]), .ZN(n27) );
  OAI211_X1 U45 ( .C1(n98), .C2(n31), .A(n28), .B(n27), .ZN(Y[15]) );
  AOI22_X1 U46 ( .A1(n8), .A2(IN0[14]), .B1(n2), .B2(IN0[16]), .ZN(n30) );
  AOI22_X1 U47 ( .A1(n87), .A2(IN0[13]), .B1(n1), .B2(IN0[15]), .ZN(n29) );
  OAI211_X1 U48 ( .C1(n91), .C2(n31), .A(n30), .B(n29), .ZN(Y[16]) );
  INV_X1 U49 ( .A(IN0[14]), .ZN(n36) );
  AOI22_X1 U50 ( .A1(n8), .A2(IN0[15]), .B1(n2), .B2(IN0[17]), .ZN(n33) );
  AOI22_X1 U51 ( .A1(n1), .A2(IN0[16]), .B1(n94), .B2(IN0[13]), .ZN(n32) );
  AOI22_X1 U52 ( .A1(n8), .A2(IN0[16]), .B1(n2), .B2(IN0[18]), .ZN(n35) );
  AOI22_X1 U53 ( .A1(n87), .A2(IN0[15]), .B1(n1), .B2(IN0[17]), .ZN(n34) );
  INV_X1 U54 ( .A(IN0[16]), .ZN(n43) );
  AOI22_X1 U55 ( .A1(n8), .A2(IN0[17]), .B1(n2), .B2(IN0[19]), .ZN(n38) );
  AOI22_X1 U56 ( .A1(n1), .A2(IN0[18]), .B1(n94), .B2(IN0[15]), .ZN(n37) );
  OAI211_X1 U57 ( .C1(n98), .C2(n43), .A(n38), .B(n37), .ZN(Y[19]) );
  INV_X1 U58 ( .A(IN0[0]), .ZN(n79) );
  AOI22_X1 U59 ( .A1(IN7[0]), .A2(n93), .B1(n2), .B2(IN0[1]), .ZN(n40) );
  AOI22_X1 U60 ( .A1(n87), .A2(IN6[0]), .B1(IN5[0]), .B2(n94), .ZN(n39) );
  OAI211_X1 U61 ( .C1(n7), .C2(n79), .A(n40), .B(n39), .ZN(Y[1]) );
  AOI22_X1 U62 ( .A1(n93), .A2(IN0[18]), .B1(n2), .B2(IN0[20]), .ZN(n42) );
  AOI22_X1 U63 ( .A1(n87), .A2(IN0[17]), .B1(n1), .B2(IN0[19]), .ZN(n41) );
  OAI211_X1 U64 ( .C1(n91), .C2(n43), .A(n42), .B(n41), .ZN(Y[20]) );
  INV_X1 U65 ( .A(IN0[18]), .ZN(n48) );
  AOI22_X1 U66 ( .A1(n8), .A2(IN0[19]), .B1(n2), .B2(IN0[21]), .ZN(n45) );
  AOI22_X1 U67 ( .A1(n1), .A2(IN0[20]), .B1(n94), .B2(IN0[17]), .ZN(n44) );
  OAI211_X1 U68 ( .C1(n98), .C2(n48), .A(n45), .B(n44), .ZN(Y[21]) );
  AOI22_X1 U69 ( .A1(n8), .A2(IN0[20]), .B1(n2), .B2(IN0[22]), .ZN(n47) );
  AOI22_X1 U70 ( .A1(n87), .A2(IN0[19]), .B1(n1), .B2(IN0[21]), .ZN(n46) );
  OAI211_X1 U71 ( .C1(n91), .C2(n48), .A(n47), .B(n46), .ZN(Y[22]) );
  INV_X1 U72 ( .A(IN0[20]), .ZN(n53) );
  AOI22_X1 U73 ( .A1(n8), .A2(IN0[21]), .B1(n2), .B2(IN0[23]), .ZN(n50) );
  AOI22_X1 U74 ( .A1(n1), .A2(IN0[22]), .B1(n94), .B2(IN0[19]), .ZN(n49) );
  OAI211_X1 U75 ( .C1(n98), .C2(n53), .A(n50), .B(n49), .ZN(Y[23]) );
  AOI22_X1 U76 ( .A1(n8), .A2(IN0[22]), .B1(n2), .B2(IN0[24]), .ZN(n52) );
  AOI22_X1 U77 ( .A1(n87), .A2(IN0[21]), .B1(n1), .B2(IN0[23]), .ZN(n51) );
  OAI211_X1 U78 ( .C1(n91), .C2(n53), .A(n52), .B(n51), .ZN(Y[24]) );
  INV_X1 U79 ( .A(IN0[22]), .ZN(n58) );
  AOI22_X1 U80 ( .A1(n8), .A2(IN0[23]), .B1(n2), .B2(IN0[25]), .ZN(n55) );
  AOI22_X1 U81 ( .A1(n1), .A2(IN0[24]), .B1(n94), .B2(IN0[21]), .ZN(n54) );
  OAI211_X1 U82 ( .C1(n98), .C2(n58), .A(n55), .B(n54), .ZN(Y[25]) );
  AOI22_X1 U83 ( .A1(n8), .A2(IN0[24]), .B1(n2), .B2(IN0[26]), .ZN(n57) );
  AOI22_X1 U84 ( .A1(n87), .A2(IN0[23]), .B1(n1), .B2(IN0[25]), .ZN(n56) );
  OAI211_X1 U85 ( .C1(n91), .C2(n58), .A(n57), .B(n56), .ZN(Y[26]) );
  INV_X1 U86 ( .A(IN0[24]), .ZN(n63) );
  AOI22_X1 U87 ( .A1(n8), .A2(IN0[25]), .B1(n2), .B2(IN0[27]), .ZN(n60) );
  AOI22_X1 U88 ( .A1(n1), .A2(IN0[26]), .B1(n94), .B2(IN0[23]), .ZN(n59) );
  OAI211_X1 U89 ( .C1(n98), .C2(n63), .A(n60), .B(n59), .ZN(Y[27]) );
  AOI22_X1 U90 ( .A1(n8), .A2(IN0[26]), .B1(n2), .B2(IN0[28]), .ZN(n62) );
  AOI22_X1 U91 ( .A1(n87), .A2(IN0[25]), .B1(n1), .B2(IN0[27]), .ZN(n61) );
  OAI211_X1 U92 ( .C1(n91), .C2(n63), .A(n62), .B(n61), .ZN(Y[28]) );
  INV_X1 U93 ( .A(IN0[26]), .ZN(n71) );
  AOI22_X1 U94 ( .A1(n93), .A2(IN0[27]), .B1(n2), .B2(IN0[29]), .ZN(n65) );
  AOI22_X1 U95 ( .A1(n1), .A2(IN0[28]), .B1(n94), .B2(IN0[25]), .ZN(n64) );
  OAI211_X1 U96 ( .C1(n98), .C2(n71), .A(n65), .B(n64), .ZN(Y[29]) );
  AOI22_X1 U97 ( .A1(n8), .A2(IN0[0]), .B1(n2), .B2(IN0[2]), .ZN(n67) );
  AOI22_X1 U98 ( .A1(n1), .A2(IN0[1]), .B1(n94), .B2(IN6[0]), .ZN(n66) );
  OAI211_X1 U99 ( .C1(n98), .C2(n68), .A(n67), .B(n66), .ZN(Y[2]) );
  AOI22_X1 U100 ( .A1(n93), .A2(IN0[28]), .B1(n2), .B2(IN0[30]), .ZN(n70) );
  AOI22_X1 U101 ( .A1(n87), .A2(IN0[27]), .B1(n1), .B2(IN0[29]), .ZN(n69) );
  OAI211_X1 U102 ( .C1(n91), .C2(n71), .A(n70), .B(n69), .ZN(Y[30]) );
  INV_X1 U103 ( .A(IN0[27]), .ZN(n74) );
  AOI22_X1 U104 ( .A1(n93), .A2(IN0[29]), .B1(n2), .B2(IN0[31]), .ZN(n73) );
  AOI22_X1 U105 ( .A1(n87), .A2(IN0[28]), .B1(n1), .B2(IN0[30]), .ZN(n72) );
  OAI211_X1 U106 ( .C1(n91), .C2(n74), .A(n73), .B(n72), .ZN(Y[31]) );
  AOI22_X1 U107 ( .A1(n93), .A2(IN0[1]), .B1(n2), .B2(n6), .ZN(n76) );
  AOI22_X1 U108 ( .A1(n1), .A2(IN0[2]), .B1(IN7[0]), .B2(n94), .ZN(n75) );
  OAI211_X1 U109 ( .C1(n98), .C2(n79), .A(n76), .B(n75), .ZN(Y[3]) );
  AOI22_X1 U110 ( .A1(n93), .A2(IN0[2]), .B1(n2), .B2(IN0[4]), .ZN(n78) );
  AOI22_X1 U111 ( .A1(n87), .A2(IN0[1]), .B1(n1), .B2(n6), .ZN(n77) );
  OAI211_X1 U112 ( .C1(n91), .C2(n79), .A(n78), .B(n77), .ZN(Y[4]) );
  INV_X1 U113 ( .A(IN0[2]), .ZN(n84) );
  AOI22_X1 U114 ( .A1(n93), .A2(n6), .B1(n2), .B2(IN0[5]), .ZN(n81) );
  AOI22_X1 U115 ( .A1(n1), .A2(IN0[4]), .B1(n94), .B2(IN0[1]), .ZN(n80) );
  OAI211_X1 U116 ( .C1(n98), .C2(n84), .A(n81), .B(n80), .ZN(Y[5]) );
  AOI22_X1 U117 ( .A1(n93), .A2(IN0[4]), .B1(n2), .B2(IN4[10]), .ZN(n83) );
  AOI22_X1 U118 ( .A1(n87), .A2(n6), .B1(n1), .B2(IN0[5]), .ZN(n82) );
  OAI211_X1 U119 ( .C1(n91), .C2(n84), .A(n83), .B(n82), .ZN(Y[6]) );
  INV_X1 U120 ( .A(IN0[4]), .ZN(n90) );
  AOI22_X1 U121 ( .A1(n8), .A2(IN0[5]), .B1(IN5[10]), .B2(n2), .ZN(n86) );
  AOI22_X1 U122 ( .A1(n1), .A2(IN4[10]), .B1(n94), .B2(IN0[3]), .ZN(n85) );
  OAI211_X1 U123 ( .C1(n98), .C2(n90), .A(n86), .B(n85), .ZN(Y[7]) );
  AOI22_X1 U124 ( .A1(n93), .A2(IN4[10]), .B1(n2), .B2(IN6[10]), .ZN(n89) );
  AOI22_X1 U125 ( .A1(n87), .A2(IN0[5]), .B1(IN5[10]), .B2(n1), .ZN(n88) );
  OAI211_X1 U126 ( .C1(n91), .C2(n90), .A(n89), .B(n88), .ZN(Y[8]) );
  INV_X1 U127 ( .A(IN4[10]), .ZN(n97) );
  AOI22_X1 U128 ( .A1(n8), .A2(IN5[10]), .B1(n2), .B2(IN7[10]), .ZN(n96) );
  AOI22_X1 U129 ( .A1(n1), .A2(IN6[10]), .B1(IN0[5]), .B2(n94), .ZN(n95) );
  OAI211_X1 U130 ( .C1(n98), .C2(n97), .A(n96), .B(n95), .ZN(Y[9]) );
endmodule


module MUX_2to1_N32_1 ( IN0, IN1, SEL, Y );
  input [31:0] IN0;
  input [31:0] IN1;
  output [31:0] Y;
  input SEL;
  wire   n2, n3, n4, n5;

  MUX2_X1 U1 ( .A(IN0[13]), .B(IN1[13]), .S(SEL), .Z(Y[13]) );
  BUF_X1 U2 ( .A(SEL), .Z(n5) );
  NAND2_X1 U3 ( .A1(n4), .A2(n2), .ZN(Y[7]) );
  OR2_X1 U4 ( .A1(SEL), .A2(n3), .ZN(n2) );
  INV_X1 U5 ( .A(IN0[7]), .ZN(n3) );
  NAND2_X1 U6 ( .A1(IN1[7]), .A2(SEL), .ZN(n4) );
  MUX2_X1 U7 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U8 ( .A(IN0[10]), .B(IN1[10]), .S(SEL), .Z(Y[10]) );
  MUX2_X1 U9 ( .A(IN0[11]), .B(IN1[11]), .S(SEL), .Z(Y[11]) );
  MUX2_X1 U10 ( .A(IN0[12]), .B(IN1[12]), .S(SEL), .Z(Y[12]) );
  MUX2_X1 U11 ( .A(IN0[14]), .B(IN1[14]), .S(SEL), .Z(Y[14]) );
  MUX2_X1 U12 ( .A(IN0[15]), .B(IN1[15]), .S(SEL), .Z(Y[15]) );
  MUX2_X1 U13 ( .A(IN0[16]), .B(IN1[16]), .S(SEL), .Z(Y[16]) );
  MUX2_X1 U14 ( .A(IN0[17]), .B(IN1[17]), .S(SEL), .Z(Y[17]) );
  MUX2_X1 U15 ( .A(IN0[18]), .B(IN1[18]), .S(SEL), .Z(Y[18]) );
  MUX2_X1 U16 ( .A(IN0[19]), .B(IN1[19]), .S(SEL), .Z(Y[19]) );
  MUX2_X1 U17 ( .A(IN0[1]), .B(IN1[1]), .S(n5), .Z(Y[1]) );
  MUX2_X1 U18 ( .A(IN0[20]), .B(IN1[20]), .S(n5), .Z(Y[20]) );
  MUX2_X1 U19 ( .A(IN0[21]), .B(IN1[21]), .S(n5), .Z(Y[21]) );
  MUX2_X1 U20 ( .A(IN0[22]), .B(IN1[22]), .S(n5), .Z(Y[22]) );
  MUX2_X1 U21 ( .A(IN0[23]), .B(IN1[23]), .S(n5), .Z(Y[23]) );
  MUX2_X1 U22 ( .A(IN0[24]), .B(IN1[24]), .S(n5), .Z(Y[24]) );
  MUX2_X1 U23 ( .A(IN0[25]), .B(IN1[25]), .S(n5), .Z(Y[25]) );
  MUX2_X1 U24 ( .A(IN0[26]), .B(IN1[26]), .S(n5), .Z(Y[26]) );
  MUX2_X1 U25 ( .A(IN0[27]), .B(IN1[27]), .S(n5), .Z(Y[27]) );
  MUX2_X1 U26 ( .A(IN0[28]), .B(IN1[28]), .S(n5), .Z(Y[28]) );
  MUX2_X1 U27 ( .A(IN0[29]), .B(IN1[29]), .S(n5), .Z(Y[29]) );
  MUX2_X1 U28 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U29 ( .A(IN0[30]), .B(IN1[30]), .S(SEL), .Z(Y[30]) );
  MUX2_X1 U30 ( .A(IN0[31]), .B(IN1[31]), .S(SEL), .Z(Y[31]) );
  MUX2_X1 U31 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
  MUX2_X1 U32 ( .A(IN0[4]), .B(IN1[4]), .S(SEL), .Z(Y[4]) );
  MUX2_X1 U33 ( .A(IN0[5]), .B(IN1[5]), .S(SEL), .Z(Y[5]) );
  MUX2_X1 U34 ( .A(IN0[6]), .B(IN1[6]), .S(SEL), .Z(Y[6]) );
  MUX2_X1 U35 ( .A(IN0[8]), .B(IN1[8]), .S(SEL), .Z(Y[8]) );
  MUX2_X1 U36 ( .A(IN0[9]), .B(IN1[9]), .S(SEL), .Z(Y[9]) );
endmodule


module barrel_shifter_Nbit32 ( A, B, SHIFT_ROTATE, LOGIC_ARITH, LEFT_RIGHT, 
        OUTPUT );
  input [31:0] A;
  input [31:0] B;
  output [31:0] OUTPUT;
  input SHIFT_ROTATE, LOGIC_ARITH, LEFT_RIGHT;
  wire   N0, N1, \out_right[8][35] , \out_right[8][34] , \out_right[8][33] ,
         \out_right[8][32] , \out_right[8][31] , \out_right[8][30] ,
         \out_right[8][29] , \out_right[8][28] , \out_right[8][27] ,
         \out_right[8][26] , \out_right[8][25] , \out_right[8][24] ,
         \out_right[8][23] , \out_right[8][22] , \out_right[8][21] ,
         \out_right[8][20] , \out_right[8][19] , \out_right[8][18] ,
         \out_right[8][17] , \out_right[8][16] , \out_right[8][15] ,
         \out_right[8][14] , \out_right[8][13] , \out_right[8][12] ,
         \out_right[8][11] , \out_right[8][10] , \out_right[8][9] ,
         \out_right[8][8] , \out_right[8][7] , \out_right[8][6] ,
         \out_right[8][5] , \out_right[8][4] , \out_right[7][35] ,
         \out_right[7][34] , \out_right[7][33] , \out_right[7][32] ,
         \out_right[7][31] , \out_right[7][30] , \out_right[7][29] ,
         \out_right[7][28] , \out_right[7][27] , \out_right[7][26] ,
         \out_right[7][25] , \out_right[7][24] , \out_right[7][23] ,
         \out_right[7][22] , \out_right[7][21] , \out_right[7][20] ,
         \out_right[7][19] , \out_right[7][18] , \out_right[7][17] ,
         \out_right[7][16] , \out_right[7][15] , \out_right[7][14] ,
         \out_right[7][13] , \out_right[7][12] , \out_right[7][11] ,
         \out_right[7][10] , \out_right[7][9] , \out_right[7][8] ,
         \out_right[6][35] , \out_right[6][34] , \out_right[6][33] ,
         \out_right[6][32] , \out_right[6][31] , \out_right[6][30] ,
         \out_right[6][29] , \out_right[6][28] , \out_right[6][27] ,
         \out_right[6][26] , \out_right[6][25] , \out_right[6][24] ,
         \out_right[6][23] , \out_right[6][22] , \out_right[6][21] ,
         \out_right[6][20] , \out_right[6][19] , \out_right[6][18] ,
         \out_right[6][17] , \out_right[6][16] , \out_right[6][15] ,
         \out_right[6][14] , \out_right[6][13] , \out_right[6][12] ,
         \out_right[5][35] , \out_right[5][34] , \out_right[5][33] ,
         \out_right[5][32] , \out_right[5][31] , \out_right[5][30] ,
         \out_right[5][29] , \out_right[5][28] , \out_right[5][27] ,
         \out_right[5][26] , \out_right[5][25] , \out_right[5][24] ,
         \out_right[5][23] , \out_right[5][22] , \out_right[5][21] ,
         \out_right[5][20] , \out_right[5][19] , \out_right[5][18] ,
         \out_right[5][17] , \out_right[5][16] , \out_right[4][35] ,
         \out_right[4][34] , \out_right[4][33] , \out_right[4][32] ,
         \out_right[4][31] , \out_right[4][30] , \out_right[4][29] ,
         \out_right[4][28] , \out_right[4][27] , \out_right[4][26] ,
         \out_right[4][25] , \out_right[4][24] , \out_right[4][23] ,
         \out_right[4][22] , \out_right[4][21] , \out_right[4][20] ,
         \out_right[3][35] , \out_right[3][34] , \out_right[3][33] ,
         \out_right[3][32] , \out_right[3][31] , \out_right[3][30] ,
         \out_right[3][29] , \out_right[3][28] , \out_right[3][27] ,
         \out_right[3][26] , \out_right[3][25] , \out_right[3][24] ,
         \out_right[2][35] , \out_right[2][34] , \out_right[2][33] ,
         \out_right[2][32] , \out_right[2][31] , \out_right[2][30] ,
         \out_right[2][29] , \out_right[2][28] , \out_right[1][35] ,
         \out_right[1][34] , \out_right[1][33] , \out_right[1][32] ,
         \out_first_stage[8][35] , \out_first_stage[8][34] ,
         \out_first_stage[8][33] , \out_first_stage[8][32] ,
         \out_first_stage[8][31] , \out_first_stage[8][30] ,
         \out_first_stage[8][29] , \out_first_stage[8][28] ,
         \out_first_stage[8][27] , \out_first_stage[8][26] ,
         \out_first_stage[8][25] , \out_first_stage[8][24] ,
         \out_first_stage[8][23] , \out_first_stage[8][22] ,
         \out_first_stage[8][21] , \out_first_stage[8][20] ,
         \out_first_stage[8][19] , \out_first_stage[8][18] ,
         \out_first_stage[8][17] , \out_first_stage[8][16] ,
         \out_first_stage[8][15] , \out_first_stage[8][14] ,
         \out_first_stage[8][13] , \out_first_stage[8][12] ,
         \out_first_stage[8][11] , \out_first_stage[8][10] ,
         \out_first_stage[8][9] , \out_first_stage[8][8] ,
         \out_first_stage[8][7] , \out_first_stage[8][6] ,
         \out_first_stage[8][5] , \out_first_stage[8][4] ,
         \out_first_stage[8][3] , \out_first_stage[8][2] ,
         \out_first_stage[8][1] , \out_first_stage[8][0] ,
         \out_first_stage[7][35] , \out_first_stage[7][34] ,
         \out_first_stage[7][33] , \out_first_stage[7][32] ,
         \out_first_stage[7][31] , \out_first_stage[7][30] ,
         \out_first_stage[7][29] , \out_first_stage[7][28] ,
         \out_first_stage[7][27] , \out_first_stage[7][26] ,
         \out_first_stage[7][25] , \out_first_stage[7][24] ,
         \out_first_stage[7][23] , \out_first_stage[7][22] ,
         \out_first_stage[7][21] , \out_first_stage[7][20] ,
         \out_first_stage[7][19] , \out_first_stage[7][18] ,
         \out_first_stage[7][17] , \out_first_stage[7][16] ,
         \out_first_stage[7][15] , \out_first_stage[7][14] ,
         \out_first_stage[7][13] , \out_first_stage[7][12] ,
         \out_first_stage[7][11] , \out_first_stage[7][10] ,
         \out_first_stage[7][9] , \out_first_stage[7][8] ,
         \out_first_stage[7][7] , \out_first_stage[7][6] ,
         \out_first_stage[7][5] , \out_first_stage[7][4] ,
         \out_first_stage[7][3] , \out_first_stage[7][2] ,
         \out_first_stage[7][1] , \out_first_stage[7][0] ,
         \out_first_stage[6][35] , \out_first_stage[6][34] ,
         \out_first_stage[6][33] , \out_first_stage[6][32] ,
         \out_first_stage[6][31] , \out_first_stage[6][30] ,
         \out_first_stage[6][29] , \out_first_stage[6][28] ,
         \out_first_stage[6][27] , \out_first_stage[6][26] ,
         \out_first_stage[6][25] , \out_first_stage[6][24] ,
         \out_first_stage[6][23] , \out_first_stage[6][22] ,
         \out_first_stage[6][21] , \out_first_stage[6][20] ,
         \out_first_stage[6][19] , \out_first_stage[6][18] ,
         \out_first_stage[6][17] , \out_first_stage[6][16] ,
         \out_first_stage[6][15] , \out_first_stage[6][14] ,
         \out_first_stage[6][13] , \out_first_stage[6][12] ,
         \out_first_stage[6][11] , \out_first_stage[6][10] ,
         \out_first_stage[6][9] , \out_first_stage[6][8] ,
         \out_first_stage[6][7] , \out_first_stage[6][6] ,
         \out_first_stage[6][5] , \out_first_stage[6][4] ,
         \out_first_stage[6][3] , \out_first_stage[6][2] ,
         \out_first_stage[6][1] , \out_first_stage[6][0] ,
         \out_first_stage[5][35] , \out_first_stage[5][34] ,
         \out_first_stage[5][33] , \out_first_stage[5][32] ,
         \out_first_stage[5][31] , \out_first_stage[5][30] ,
         \out_first_stage[5][29] , \out_first_stage[5][28] ,
         \out_first_stage[5][27] , \out_first_stage[5][26] ,
         \out_first_stage[5][25] , \out_first_stage[5][24] ,
         \out_first_stage[5][23] , \out_first_stage[5][22] ,
         \out_first_stage[5][21] , \out_first_stage[5][20] ,
         \out_first_stage[5][19] , \out_first_stage[5][18] ,
         \out_first_stage[5][17] , \out_first_stage[5][16] ,
         \out_first_stage[5][15] , \out_first_stage[5][14] ,
         \out_first_stage[5][13] , \out_first_stage[5][12] ,
         \out_first_stage[5][11] , \out_first_stage[5][10] ,
         \out_first_stage[5][9] , \out_first_stage[5][8] ,
         \out_first_stage[5][7] , \out_first_stage[5][6] ,
         \out_first_stage[5][5] , \out_first_stage[5][4] ,
         \out_first_stage[5][3] , \out_first_stage[5][2] ,
         \out_first_stage[5][1] , \out_first_stage[5][0] ,
         \out_first_stage[4][35] , \out_first_stage[4][34] ,
         \out_first_stage[4][33] , \out_first_stage[4][32] ,
         \out_first_stage[4][31] , \out_first_stage[4][30] ,
         \out_first_stage[4][29] , \out_first_stage[4][28] ,
         \out_first_stage[4][27] , \out_first_stage[4][26] ,
         \out_first_stage[4][25] , \out_first_stage[4][24] ,
         \out_first_stage[4][23] , \out_first_stage[4][22] ,
         \out_first_stage[4][21] , \out_first_stage[4][20] ,
         \out_first_stage[4][19] , \out_first_stage[4][18] ,
         \out_first_stage[4][17] , \out_first_stage[4][16] ,
         \out_first_stage[4][15] , \out_first_stage[4][14] ,
         \out_first_stage[4][13] , \out_first_stage[4][12] ,
         \out_first_stage[4][11] , \out_first_stage[4][10] ,
         \out_first_stage[4][9] , \out_first_stage[4][8] ,
         \out_first_stage[4][7] , \out_first_stage[4][6] ,
         \out_first_stage[4][5] , \out_first_stage[4][4] ,
         \out_first_stage[4][3] , \out_first_stage[4][2] ,
         \out_first_stage[4][1] , \out_first_stage[4][0] ,
         \out_first_stage[3][35] , \out_first_stage[3][34] ,
         \out_first_stage[3][33] , \out_first_stage[3][32] ,
         \out_first_stage[3][31] , \out_first_stage[3][30] ,
         \out_first_stage[3][29] , \out_first_stage[3][28] ,
         \out_first_stage[3][27] , \out_first_stage[3][26] ,
         \out_first_stage[3][25] , \out_first_stage[3][24] ,
         \out_first_stage[3][23] , \out_first_stage[3][22] ,
         \out_first_stage[3][21] , \out_first_stage[3][20] ,
         \out_first_stage[3][19] , \out_first_stage[3][18] ,
         \out_first_stage[3][17] , \out_first_stage[3][16] ,
         \out_first_stage[3][15] , \out_first_stage[3][14] ,
         \out_first_stage[3][13] , \out_first_stage[3][12] ,
         \out_first_stage[3][11] , \out_first_stage[3][10] ,
         \out_first_stage[3][9] , \out_first_stage[3][8] ,
         \out_first_stage[3][7] , \out_first_stage[3][6] ,
         \out_first_stage[3][5] , \out_first_stage[3][4] ,
         \out_first_stage[3][3] , \out_first_stage[3][2] ,
         \out_first_stage[3][1] , \out_first_stage[3][0] ,
         \out_first_stage[2][35] , \out_first_stage[2][34] ,
         \out_first_stage[2][33] , \out_first_stage[2][32] ,
         \out_first_stage[2][31] , \out_first_stage[2][30] ,
         \out_first_stage[2][29] , \out_first_stage[2][28] ,
         \out_first_stage[2][27] , \out_first_stage[2][26] ,
         \out_first_stage[2][25] , \out_first_stage[2][24] ,
         \out_first_stage[2][23] , \out_first_stage[2][22] ,
         \out_first_stage[2][21] , \out_first_stage[2][20] ,
         \out_first_stage[2][19] , \out_first_stage[2][18] ,
         \out_first_stage[2][17] , \out_first_stage[2][16] ,
         \out_first_stage[2][15] , \out_first_stage[2][14] ,
         \out_first_stage[2][13] , \out_first_stage[2][12] ,
         \out_first_stage[2][11] , \out_first_stage[2][10] ,
         \out_first_stage[2][9] , \out_first_stage[2][8] ,
         \out_first_stage[2][7] , \out_first_stage[2][6] ,
         \out_first_stage[2][5] , \out_first_stage[2][4] ,
         \out_first_stage[2][3] , \out_first_stage[2][2] ,
         \out_first_stage[2][1] , \out_first_stage[2][0] ,
         \out_first_stage[1][35] , \out_first_stage[1][34] ,
         \out_first_stage[1][33] , \out_first_stage[1][32] ,
         \out_first_stage[1][31] , \out_first_stage[1][30] ,
         \out_first_stage[1][29] , \out_first_stage[1][28] ,
         \out_first_stage[1][27] , \out_first_stage[1][26] ,
         \out_first_stage[1][25] , \out_first_stage[1][24] ,
         \out_first_stage[1][23] , \out_first_stage[1][22] ,
         \out_first_stage[1][21] , \out_first_stage[1][20] ,
         \out_first_stage[1][19] , \out_first_stage[1][18] ,
         \out_first_stage[1][17] , \out_first_stage[1][16] ,
         \out_first_stage[1][15] , \out_first_stage[1][14] ,
         \out_first_stage[1][13] , \out_first_stage[1][12] ,
         \out_first_stage[1][11] , \out_first_stage[1][10] ,
         \out_first_stage[1][9] , \out_first_stage[1][8] ,
         \out_first_stage[1][7] , \out_first_stage[1][6] ,
         \out_first_stage[1][5] , \out_first_stage[1][4] ,
         \out_first_stage[1][3] , \out_first_stage[1][2] ,
         \out_first_stage[1][1] , \out_first_stage[1][0] , n9, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320;
  wire   [31:0] out_control;
  wire   [4:0] shift_pos;
  wire   [31:0] fill_vector_left;
  wire   [31:0] fill_vector_right;
  wire   [35:0] out_second_stage;
  wire   [31:0] out_barrel;

  MUX_2to1_N32_4 mux_shift_rotate_left ( .IN0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .IN1(A), .SEL(SHIFT_ROTATE), .Y(fill_vector_left)
         );
  MUX_2to1_N32_3 mux_shift_rotate_right ( .IN0({A[31], A[31], A[31], A[31], 
        A[31], A[31], A[31], A[31], A[31], A[31], A[31], A[31], A[31], A[31], 
        A[31], A[31], A[31], A[31], A[31], A[31], A[31], A[31], A[31], A[31], 
        A[31], A[31], A[31], A[31], A[31], A[31], A[31], A[31]}), .IN1({1'b0, 
        A[30:0]}), .SEL(SHIFT_ROTATE), .Y(fill_vector_right) );
  MUX_2to1_N4_0 right_MUX2to1_1 ( .IN0({1'b0, 1'b0, 1'b0, 1'b0}), .IN1(
        fill_vector_right[3:0]), .SEL(n311), .Y({\out_right[1][35] , 
        \out_right[1][34] , \out_right[1][33] , \out_right[1][32] }) );
  MUX_2to1_N8 right_MUX2to1_2 ( .IN0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .IN1(fill_vector_right[7:0]), .SEL(n311), .Y({
        \out_right[2][35] , \out_right[2][34] , \out_right[2][33] , 
        \out_right[2][32] , \out_right[2][31] , \out_right[2][30] , 
        \out_right[2][29] , \out_right[2][28] }) );
  MUX_2to1_N12 right_MUX2to1_3 ( .IN0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN1(fill_vector_right[11:0]), 
        .SEL(n311), .Y({\out_right[3][35] , \out_right[3][34] , 
        \out_right[3][33] , \out_right[3][32] , \out_right[3][31] , 
        \out_right[3][30] , \out_right[3][29] , \out_right[3][28] , 
        \out_right[3][27] , \out_right[3][26] , \out_right[3][25] , 
        \out_right[3][24] }) );
  MUX_2to1_N16 right_MUX2to1_4 ( .IN0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN1(
        fill_vector_right[15:0]), .SEL(n311), .Y({\out_right[4][35] , 
        \out_right[4][34] , \out_right[4][33] , \out_right[4][32] , 
        \out_right[4][31] , \out_right[4][30] , \out_right[4][29] , 
        \out_right[4][28] , \out_right[4][27] , \out_right[4][26] , 
        \out_right[4][25] , \out_right[4][24] , \out_right[4][23] , 
        \out_right[4][22] , \out_right[4][21] , \out_right[4][20] }) );
  MUX_2to1_N20 right_MUX2to1_5 ( .IN0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .IN1(fill_vector_right[19:0]), .SEL(n311), .Y({
        \out_right[5][35] , \out_right[5][34] , \out_right[5][33] , 
        \out_right[5][32] , \out_right[5][31] , \out_right[5][30] , 
        \out_right[5][29] , \out_right[5][28] , \out_right[5][27] , 
        \out_right[5][26] , \out_right[5][25] , \out_right[5][24] , 
        \out_right[5][23] , \out_right[5][22] , \out_right[5][21] , 
        \out_right[5][20] , \out_right[5][19] , \out_right[5][18] , 
        \out_right[5][17] , \out_right[5][16] }) );
  MUX_2to1_N24 right_MUX2to1_6 ( .IN0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN1(fill_vector_right[23:0]), 
        .SEL(LOGIC_ARITH), .Y({\out_right[6][35] , \out_right[6][34] , 
        \out_right[6][33] , \out_right[6][32] , \out_right[6][31] , 
        \out_right[6][30] , \out_right[6][29] , \out_right[6][28] , 
        \out_right[6][27] , \out_right[6][26] , \out_right[6][25] , 
        \out_right[6][24] , \out_right[6][23] , \out_right[6][22] , 
        \out_right[6][21] , \out_right[6][20] , \out_right[6][19] , 
        \out_right[6][18] , \out_right[6][17] , \out_right[6][16] , 
        \out_right[6][15] , \out_right[6][14] , \out_right[6][13] , 
        \out_right[6][12] }) );
  MUX_2to1_N28 right_MUX2to1_7 ( .IN0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN1(
        fill_vector_right[27:0]), .SEL(LOGIC_ARITH), .Y({\out_right[7][35] , 
        \out_right[7][34] , \out_right[7][33] , \out_right[7][32] , 
        \out_right[7][31] , \out_right[7][30] , \out_right[7][29] , 
        \out_right[7][28] , \out_right[7][27] , \out_right[7][26] , 
        \out_right[7][25] , \out_right[7][24] , \out_right[7][23] , 
        \out_right[7][22] , \out_right[7][21] , \out_right[7][20] , 
        \out_right[7][19] , \out_right[7][18] , \out_right[7][17] , 
        \out_right[7][16] , \out_right[7][15] , \out_right[7][14] , 
        \out_right[7][13] , \out_right[7][12] , \out_right[7][11] , 
        \out_right[7][10] , \out_right[7][9] , \out_right[7][8] }) );
  MUX_2to1_N32_2 right_MUX2to1_8 ( .IN0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .IN1(fill_vector_right), .SEL(n311), .Y({
        \out_right[8][35] , \out_right[8][34] , \out_right[8][33] , 
        \out_right[8][32] , \out_right[8][31] , \out_right[8][30] , 
        \out_right[8][29] , \out_right[8][28] , \out_right[8][27] , 
        \out_right[8][26] , \out_right[8][25] , \out_right[8][24] , 
        \out_right[8][23] , \out_right[8][22] , \out_right[8][21] , 
        \out_right[8][20] , \out_right[8][19] , \out_right[8][18] , 
        \out_right[8][17] , \out_right[8][16] , \out_right[8][15] , 
        \out_right[8][14] , \out_right[8][13] , \out_right[8][12] , 
        \out_right[8][11] , \out_right[8][10] , \out_right[8][9] , 
        \out_right[8][8] , \out_right[8][7] , \out_right[8][6] , 
        \out_right[8][5] , \out_right[8][4] }) );
  MUX_2to1_N36_0 MASK_MUX2to1_1 ( .IN0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, A[9:6], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        fill_vector_left[31:28]}), .IN1({\out_right[1][35] , 
        \out_right[1][34] , \out_right[1][33] , \out_right[1][32] , A[31:10], 
        1'b0, 1'b0, 1'b0, 1'b0, A[5:0]}), .SEL(n310), .Y({
        \out_first_stage[1][35] , \out_first_stage[1][34] , 
        \out_first_stage[1][33] , \out_first_stage[1][32] , 
        \out_first_stage[1][31] , \out_first_stage[1][30] , 
        \out_first_stage[1][29] , \out_first_stage[1][28] , 
        \out_first_stage[1][27] , \out_first_stage[1][26] , 
        \out_first_stage[1][25] , \out_first_stage[1][24] , 
        \out_first_stage[1][23] , \out_first_stage[1][22] , 
        \out_first_stage[1][21] , \out_first_stage[1][20] , 
        \out_first_stage[1][19] , \out_first_stage[1][18] , 
        \out_first_stage[1][17] , \out_first_stage[1][16] , 
        \out_first_stage[1][15] , \out_first_stage[1][14] , 
        \out_first_stage[1][13] , \out_first_stage[1][12] , 
        \out_first_stage[1][11] , \out_first_stage[1][10] , 
        \out_first_stage[1][9] , \out_first_stage[1][8] , 
        \out_first_stage[1][7] , \out_first_stage[1][6] , 
        \out_first_stage[1][5] , \out_first_stage[1][4] , 
        \out_first_stage[1][3] , \out_first_stage[1][2] , 
        \out_first_stage[1][1] , \out_first_stage[1][0] }) );
  MUX_2to1_N36_7 MASK_MUX2to1_2 ( .IN0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, A[13:5], 1'b0, A[3:0], 
        fill_vector_left[31:24]}), .IN1({\out_right[2][35] , 
        \out_right[2][34] , \out_right[2][33] , \out_right[2][32] , 
        \out_right[2][31] , \out_right[2][30] , \out_right[2][29] , 
        \out_right[2][28] , A[31:14], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, A[4]}), .SEL(n310), .Y({\out_first_stage[2][35] , 
        \out_first_stage[2][34] , \out_first_stage[2][33] , 
        \out_first_stage[2][32] , \out_first_stage[2][31] , 
        \out_first_stage[2][30] , \out_first_stage[2][29] , 
        \out_first_stage[2][28] , \out_first_stage[2][27] , 
        \out_first_stage[2][26] , \out_first_stage[2][25] , 
        \out_first_stage[2][24] , \out_first_stage[2][23] , 
        \out_first_stage[2][22] , \out_first_stage[2][21] , 
        \out_first_stage[2][20] , \out_first_stage[2][19] , 
        \out_first_stage[2][18] , \out_first_stage[2][17] , 
        \out_first_stage[2][16] , \out_first_stage[2][15] , 
        \out_first_stage[2][14] , \out_first_stage[2][13] , 
        \out_first_stage[2][12] , \out_first_stage[2][11] , 
        \out_first_stage[2][10] , \out_first_stage[2][9] , 
        \out_first_stage[2][8] , \out_first_stage[2][7] , 
        \out_first_stage[2][6] , \out_first_stage[2][5] , 
        \out_first_stage[2][4] , \out_first_stage[2][3] , 
        \out_first_stage[2][2] , \out_first_stage[2][1] , 
        \out_first_stage[2][0] }) );
  MUX_2to1_N36_6 MASK_MUX2to1_3 ( .IN0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        A[17:10], 1'b0, 1'b0, A[7:0], fill_vector_left[31:20]}), .IN1({
        \out_right[3][35] , \out_right[3][34] , \out_right[3][33] , 
        \out_right[3][32] , \out_right[3][31] , \out_right[3][30] , 
        \out_right[3][29] , \out_right[3][28] , \out_right[3][27] , 
        \out_right[3][26] , \out_right[3][25] , \out_right[3][24] , A[31:18], 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, A[9:8]}), .SEL(n310), 
        .Y({\out_first_stage[3][35] , \out_first_stage[3][34] , 
        \out_first_stage[3][33] , \out_first_stage[3][32] , 
        \out_first_stage[3][31] , \out_first_stage[3][30] , 
        \out_first_stage[3][29] , \out_first_stage[3][28] , 
        \out_first_stage[3][27] , \out_first_stage[3][26] , 
        \out_first_stage[3][25] , \out_first_stage[3][24] , 
        \out_first_stage[3][23] , \out_first_stage[3][22] , 
        \out_first_stage[3][21] , \out_first_stage[3][20] , 
        \out_first_stage[3][19] , \out_first_stage[3][18] , 
        \out_first_stage[3][17] , \out_first_stage[3][16] , 
        \out_first_stage[3][15] , \out_first_stage[3][14] , 
        \out_first_stage[3][13] , \out_first_stage[3][12] , 
        \out_first_stage[3][11] , \out_first_stage[3][10] , 
        \out_first_stage[3][9] , \out_first_stage[3][8] , 
        \out_first_stage[3][7] , \out_first_stage[3][6] , 
        \out_first_stage[3][5] , \out_first_stage[3][4] , 
        \out_first_stage[3][3] , \out_first_stage[3][2] , 
        \out_first_stage[3][1] , \out_first_stage[3][0] }) );
  MUX_2to1_N36_5 MASK_MUX2to1_4 ( .IN0({A[19:15], 1'b0, 1'b0, 1'b0, A[11:0], 
        fill_vector_left[31:16]}), .IN1({\out_right[4][35] , 
        \out_right[4][34] , \out_right[4][33] , \out_right[4][32] , 
        \out_right[4][31] , \out_right[4][30] , \out_right[4][29] , 
        \out_right[4][28] , \out_right[4][27] , \out_right[4][26] , 
        \out_right[4][25] , \out_right[4][24] , \out_right[4][23] , 
        \out_right[4][22] , \out_right[4][21] , \out_right[4][20] , A[31:20], 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, A[14:12]}), .SEL(n310), .Y({
        \out_first_stage[4][35] , \out_first_stage[4][34] , 
        \out_first_stage[4][33] , \out_first_stage[4][32] , 
        \out_first_stage[4][31] , \out_first_stage[4][30] , 
        \out_first_stage[4][29] , \out_first_stage[4][28] , 
        \out_first_stage[4][27] , \out_first_stage[4][26] , 
        \out_first_stage[4][25] , \out_first_stage[4][24] , 
        \out_first_stage[4][23] , \out_first_stage[4][22] , 
        \out_first_stage[4][21] , \out_first_stage[4][20] , 
        \out_first_stage[4][19] , \out_first_stage[4][18] , 
        \out_first_stage[4][17] , \out_first_stage[4][16] , 
        \out_first_stage[4][15] , \out_first_stage[4][14] , 
        \out_first_stage[4][13] , \out_first_stage[4][12] , 
        \out_first_stage[4][11] , \out_first_stage[4][10] , 
        \out_first_stage[4][9] , \out_first_stage[4][8] , 
        \out_first_stage[4][7] , \out_first_stage[4][6] , 
        \out_first_stage[4][5] , \out_first_stage[4][4] , 
        \out_first_stage[4][3] , \out_first_stage[4][2] , 
        \out_first_stage[4][1] , \out_first_stage[4][0] }) );
  MUX_2to1_N36_4 MASK_MUX2to1_5 ( .IN0({A[15:0], fill_vector_left[31:12]}), 
        .IN1({\out_right[5][35] , \out_right[5][34] , \out_right[5][33] , 
        \out_right[5][32] , \out_right[5][31] , \out_right[5][30] , 
        \out_right[5][29] , \out_right[5][28] , \out_right[5][27] , 
        \out_right[5][26] , \out_right[5][25] , \out_right[5][24] , 
        \out_right[5][23] , \out_right[5][22] , \out_right[5][21] , 
        \out_right[5][20] , \out_right[5][19] , \out_right[5][18] , 
        \out_right[5][17] , \out_right[5][16] , A[31:16]}), .SEL(n310), .Y({
        \out_first_stage[5][35] , \out_first_stage[5][34] , 
        \out_first_stage[5][33] , \out_first_stage[5][32] , 
        \out_first_stage[5][31] , \out_first_stage[5][30] , 
        \out_first_stage[5][29] , \out_first_stage[5][28] , 
        \out_first_stage[5][27] , \out_first_stage[5][26] , 
        \out_first_stage[5][25] , \out_first_stage[5][24] , 
        \out_first_stage[5][23] , \out_first_stage[5][22] , 
        \out_first_stage[5][21] , \out_first_stage[5][20] , 
        \out_first_stage[5][19] , \out_first_stage[5][18] , 
        \out_first_stage[5][17] , \out_first_stage[5][16] , 
        \out_first_stage[5][15] , \out_first_stage[5][14] , 
        \out_first_stage[5][13] , \out_first_stage[5][12] , 
        \out_first_stage[5][11] , \out_first_stage[5][10] , 
        \out_first_stage[5][9] , \out_first_stage[5][8] , 
        \out_first_stage[5][7] , \out_first_stage[5][6] , 
        \out_first_stage[5][5] , \out_first_stage[5][4] , 
        \out_first_stage[5][3] , \out_first_stage[5][2] , 
        \out_first_stage[5][1] , \out_first_stage[5][0] }) );
  MUX_2to1_N36_3 MASK_MUX2to1_6 ( .IN0({A[11:0], fill_vector_left[31:8]}), 
        .IN1({\out_right[6][35] , \out_right[6][34] , \out_right[6][33] , 
        \out_right[6][32] , \out_right[6][31] , \out_right[6][30] , 
        \out_right[6][29] , \out_right[6][28] , \out_right[6][27] , 
        \out_right[6][26] , \out_right[6][25] , \out_right[6][24] , 
        \out_right[6][23] , \out_right[6][22] , \out_right[6][21] , 
        \out_right[6][20] , \out_right[6][19] , \out_right[6][18] , 
        \out_right[6][17] , \out_right[6][16] , \out_right[6][15] , 
        \out_right[6][14] , \out_right[6][13] , \out_right[6][12] , A[31:20]}), 
        .SEL(n310), .Y({\out_first_stage[6][35] , \out_first_stage[6][34] , 
        \out_first_stage[6][33] , \out_first_stage[6][32] , 
        \out_first_stage[6][31] , \out_first_stage[6][30] , 
        \out_first_stage[6][29] , \out_first_stage[6][28] , 
        \out_first_stage[6][27] , \out_first_stage[6][26] , 
        \out_first_stage[6][25] , \out_first_stage[6][24] , 
        \out_first_stage[6][23] , \out_first_stage[6][22] , 
        \out_first_stage[6][21] , \out_first_stage[6][20] , 
        \out_first_stage[6][19] , \out_first_stage[6][18] , 
        \out_first_stage[6][17] , \out_first_stage[6][16] , 
        \out_first_stage[6][15] , \out_first_stage[6][14] , 
        \out_first_stage[6][13] , \out_first_stage[6][12] , 
        \out_first_stage[6][11] , \out_first_stage[6][10] , 
        \out_first_stage[6][9] , \out_first_stage[6][8] , 
        \out_first_stage[6][7] , \out_first_stage[6][6] , 
        \out_first_stage[6][5] , \out_first_stage[6][4] , 
        \out_first_stage[6][3] , \out_first_stage[6][2] , 
        \out_first_stage[6][1] , \out_first_stage[6][0] }) );
  MUX_2to1_N36_2 MASK_MUX2to1_7 ( .IN0({A[7:0], fill_vector_left[31:4]}), 
        .IN1({\out_right[7][35] , \out_right[7][34] , \out_right[7][33] , 
        \out_right[7][32] , \out_right[7][31] , \out_right[7][30] , 
        \out_right[7][29] , \out_right[7][28] , \out_right[7][27] , 
        \out_right[7][26] , \out_right[7][25] , \out_right[7][24] , 
        \out_right[7][23] , \out_right[7][22] , \out_right[7][21] , 
        \out_right[7][20] , \out_right[7][19] , \out_right[7][18] , 
        \out_right[7][17] , \out_right[7][16] , \out_right[7][15] , 
        \out_right[7][14] , \out_right[7][13] , \out_right[7][12] , 
        \out_right[7][11] , \out_right[7][10] , \out_right[7][9] , 
        \out_right[7][8] , A[31:24]}), .SEL(n310), .Y({
        \out_first_stage[7][35] , \out_first_stage[7][34] , 
        \out_first_stage[7][33] , \out_first_stage[7][32] , 
        \out_first_stage[7][31] , \out_first_stage[7][30] , 
        \out_first_stage[7][29] , \out_first_stage[7][28] , 
        \out_first_stage[7][27] , \out_first_stage[7][26] , 
        \out_first_stage[7][25] , \out_first_stage[7][24] , 
        \out_first_stage[7][23] , \out_first_stage[7][22] , 
        \out_first_stage[7][21] , \out_first_stage[7][20] , 
        \out_first_stage[7][19] , \out_first_stage[7][18] , 
        \out_first_stage[7][17] , \out_first_stage[7][16] , 
        \out_first_stage[7][15] , \out_first_stage[7][14] , 
        \out_first_stage[7][13] , \out_first_stage[7][12] , 
        \out_first_stage[7][11] , \out_first_stage[7][10] , 
        \out_first_stage[7][9] , \out_first_stage[7][8] , 
        \out_first_stage[7][7] , \out_first_stage[7][6] , 
        \out_first_stage[7][5] , \out_first_stage[7][4] , 
        \out_first_stage[7][3] , \out_first_stage[7][2] , 
        \out_first_stage[7][1] , \out_first_stage[7][0] }) );
  MUX_2to1_N36_1 MASK_MUX2to1_8 ( .IN0({A[3:0], fill_vector_left}), .IN1({
        \out_right[8][35] , \out_right[8][34] , \out_right[8][33] , 
        \out_right[8][32] , \out_right[8][31] , \out_right[8][30] , 
        \out_right[8][29] , \out_right[8][28] , \out_right[8][27] , 
        \out_right[8][26] , \out_right[8][25] , \out_right[8][24] , 
        \out_right[8][23] , \out_right[8][22] , \out_right[8][21] , 
        \out_right[8][20] , \out_right[8][19] , \out_right[8][18] , 
        \out_right[8][17] , \out_right[8][16] , \out_right[8][15] , 
        \out_right[8][14] , \out_right[8][13] , \out_right[8][12] , 
        \out_right[8][11] , \out_right[8][10] , \out_right[8][9] , 
        \out_right[8][8] , \out_right[8][7] , \out_right[8][6] , 
        \out_right[8][5] , \out_right[8][4] , A[31:28]}), .SEL(n310), .Y({
        \out_first_stage[8][35] , \out_first_stage[8][34] , 
        \out_first_stage[8][33] , \out_first_stage[8][32] , 
        \out_first_stage[8][31] , \out_first_stage[8][30] , 
        \out_first_stage[8][29] , \out_first_stage[8][28] , 
        \out_first_stage[8][27] , \out_first_stage[8][26] , 
        \out_first_stage[8][25] , \out_first_stage[8][24] , 
        \out_first_stage[8][23] , \out_first_stage[8][22] , 
        \out_first_stage[8][21] , \out_first_stage[8][20] , 
        \out_first_stage[8][19] , \out_first_stage[8][18] , 
        \out_first_stage[8][17] , \out_first_stage[8][16] , 
        \out_first_stage[8][15] , \out_first_stage[8][14] , 
        \out_first_stage[8][13] , \out_first_stage[8][12] , 
        \out_first_stage[8][11] , \out_first_stage[8][10] , 
        \out_first_stage[8][9] , \out_first_stage[8][8] , 
        \out_first_stage[8][7] , \out_first_stage[8][6] , 
        \out_first_stage[8][5] , \out_first_stage[8][4] , 
        \out_first_stage[8][3] , \out_first_stage[8][2] , 
        \out_first_stage[8][1] , \out_first_stage[8][0] }) );
  MUX_8to1_N36 mux_second_stage ( .IN0({\out_first_stage[1][35] , 
        \out_first_stage[1][34] , \out_first_stage[1][33] , 
        \out_first_stage[1][32] , \out_first_stage[1][31] , 
        \out_first_stage[1][30] , \out_first_stage[1][29] , 
        \out_first_stage[1][28] , \out_first_stage[1][27] , 
        \out_first_stage[1][26] , \out_first_stage[1][25] , 
        \out_first_stage[1][24] , \out_first_stage[1][23] , 
        \out_first_stage[1][22] , \out_first_stage[1][21] , 
        \out_first_stage[1][20] , \out_first_stage[1][19] , 
        \out_first_stage[1][18] , \out_first_stage[1][17] , 
        \out_first_stage[1][16] , \out_first_stage[1][15] , 
        \out_first_stage[1][14] , \out_first_stage[1][13] , 
        \out_first_stage[1][12] , \out_first_stage[1][11] , 
        \out_first_stage[1][10] , \out_first_stage[1][9] , 
        \out_first_stage[1][8] , \out_first_stage[1][7] , 
        \out_first_stage[1][6] , \out_first_stage[1][5] , 
        \out_first_stage[1][4] , \out_first_stage[1][3] , 
        \out_first_stage[1][2] , \out_first_stage[1][1] , 
        \out_first_stage[1][0] }), .IN1({\out_first_stage[2][35] , 
        \out_first_stage[2][34] , \out_first_stage[2][33] , 
        \out_first_stage[2][32] , \out_first_stage[2][31] , 
        \out_first_stage[2][30] , \out_first_stage[2][29] , 
        \out_first_stage[2][28] , \out_first_stage[2][27] , 
        \out_first_stage[2][26] , \out_first_stage[2][25] , 
        \out_first_stage[2][24] , \out_first_stage[2][23] , 
        \out_first_stage[2][22] , \out_first_stage[2][21] , 
        \out_first_stage[2][20] , \out_first_stage[2][19] , 
        \out_first_stage[2][18] , \out_first_stage[2][17] , 
        \out_first_stage[2][16] , \out_first_stage[2][15] , 
        \out_first_stage[2][14] , \out_first_stage[2][13] , 
        \out_first_stage[2][12] , \out_first_stage[2][11] , 
        \out_first_stage[2][10] , \out_first_stage[2][9] , 
        \out_first_stage[2][8] , \out_first_stage[2][7] , 
        \out_first_stage[2][6] , \out_first_stage[2][5] , 
        \out_first_stage[2][4] , \out_first_stage[2][3] , 
        \out_first_stage[2][2] , \out_first_stage[2][1] , 
        \out_first_stage[2][0] }), .IN2({\out_first_stage[3][35] , 
        \out_first_stage[3][34] , \out_first_stage[3][33] , 
        \out_first_stage[3][32] , \out_first_stage[3][31] , 
        \out_first_stage[3][30] , \out_first_stage[3][29] , 
        \out_first_stage[3][28] , \out_first_stage[3][27] , 
        \out_first_stage[3][26] , \out_first_stage[3][25] , 
        \out_first_stage[3][24] , \out_first_stage[3][23] , 
        \out_first_stage[3][22] , \out_first_stage[3][21] , 
        \out_first_stage[3][20] , \out_first_stage[3][19] , 
        \out_first_stage[3][18] , \out_first_stage[3][17] , 
        \out_first_stage[3][16] , \out_first_stage[3][15] , 
        \out_first_stage[3][14] , \out_first_stage[3][13] , 
        \out_first_stage[3][12] , \out_first_stage[3][11] , 
        \out_first_stage[3][10] , \out_first_stage[3][9] , 
        \out_first_stage[3][8] , \out_first_stage[3][7] , 
        \out_first_stage[3][6] , \out_first_stage[3][5] , 
        \out_first_stage[3][4] , \out_first_stage[3][3] , 
        \out_first_stage[3][2] , \out_first_stage[3][1] , 
        \out_first_stage[3][0] }), .IN3({\out_first_stage[4][35] , 
        \out_first_stage[4][34] , \out_first_stage[4][33] , 
        \out_first_stage[4][32] , \out_first_stage[4][31] , 
        \out_first_stage[4][30] , \out_first_stage[4][29] , 
        \out_first_stage[4][28] , \out_first_stage[4][27] , 
        \out_first_stage[4][26] , \out_first_stage[4][25] , 
        \out_first_stage[4][24] , \out_first_stage[4][23] , 
        \out_first_stage[4][22] , \out_first_stage[4][21] , 
        \out_first_stage[4][20] , \out_first_stage[4][19] , 
        \out_first_stage[4][18] , \out_first_stage[4][17] , 
        \out_first_stage[4][16] , \out_first_stage[4][15] , 
        \out_first_stage[4][14] , \out_first_stage[4][13] , 
        \out_first_stage[4][12] , \out_first_stage[4][11] , 
        \out_first_stage[4][10] , \out_first_stage[4][9] , 
        \out_first_stage[4][8] , \out_first_stage[4][7] , 
        \out_first_stage[4][6] , \out_first_stage[4][5] , 
        \out_first_stage[4][4] , \out_first_stage[4][3] , 
        \out_first_stage[4][2] , \out_first_stage[4][1] , 
        \out_first_stage[4][0] }), .IN4({\out_first_stage[5][35] , 
        \out_first_stage[5][34] , \out_first_stage[5][33] , 
        \out_first_stage[5][32] , \out_first_stage[5][31] , 
        \out_first_stage[5][30] , \out_first_stage[5][29] , 
        \out_first_stage[5][28] , \out_first_stage[5][27] , 
        \out_first_stage[5][26] , \out_first_stage[5][25] , 
        \out_first_stage[5][24] , \out_first_stage[5][23] , 
        \out_first_stage[5][22] , \out_first_stage[5][21] , 
        \out_first_stage[5][20] , \out_first_stage[5][19] , 
        \out_first_stage[5][18] , \out_first_stage[5][17] , 
        \out_first_stage[5][16] , \out_first_stage[5][15] , 
        \out_first_stage[5][14] , \out_first_stage[5][13] , 
        \out_first_stage[5][12] , \out_first_stage[5][11] , 
        \out_first_stage[5][10] , \out_first_stage[5][9] , 
        \out_first_stage[5][8] , \out_first_stage[5][7] , 
        \out_first_stage[5][6] , \out_first_stage[5][5] , 
        \out_first_stage[5][4] , \out_first_stage[5][3] , 
        \out_first_stage[5][2] , \out_first_stage[5][1] , 
        \out_first_stage[5][0] }), .IN5({\out_first_stage[6][35] , 
        \out_first_stage[6][34] , \out_first_stage[6][33] , 
        \out_first_stage[6][32] , \out_first_stage[6][31] , 
        \out_first_stage[6][30] , \out_first_stage[6][29] , 
        \out_first_stage[6][28] , \out_first_stage[6][27] , 
        \out_first_stage[6][26] , \out_first_stage[6][25] , 
        \out_first_stage[6][24] , \out_first_stage[6][23] , 
        \out_first_stage[6][22] , \out_first_stage[6][21] , 
        \out_first_stage[6][20] , \out_first_stage[6][19] , 
        \out_first_stage[6][18] , \out_first_stage[6][17] , 
        \out_first_stage[6][16] , \out_first_stage[6][15] , 
        \out_first_stage[6][14] , \out_first_stage[6][13] , 
        \out_first_stage[6][12] , \out_first_stage[6][11] , 
        \out_first_stage[6][10] , \out_first_stage[6][9] , 
        \out_first_stage[6][8] , \out_first_stage[6][7] , 
        \out_first_stage[6][6] , \out_first_stage[6][5] , 
        \out_first_stage[6][4] , \out_first_stage[6][3] , 
        \out_first_stage[6][2] , \out_first_stage[6][1] , 
        \out_first_stage[6][0] }), .IN6({\out_first_stage[7][35] , 
        \out_first_stage[7][34] , \out_first_stage[7][33] , 
        \out_first_stage[7][32] , \out_first_stage[7][31] , 
        \out_first_stage[7][30] , \out_first_stage[7][29] , 
        \out_first_stage[7][28] , \out_first_stage[7][27] , 
        \out_first_stage[7][26] , \out_first_stage[7][25] , 
        \out_first_stage[7][24] , \out_first_stage[7][23] , 
        \out_first_stage[7][22] , \out_first_stage[7][21] , 
        \out_first_stage[7][20] , \out_first_stage[7][19] , 
        \out_first_stage[7][18] , \out_first_stage[7][17] , 
        \out_first_stage[7][16] , \out_first_stage[7][15] , 
        \out_first_stage[7][14] , \out_first_stage[7][13] , 
        \out_first_stage[7][12] , \out_first_stage[7][11] , 
        \out_first_stage[7][10] , \out_first_stage[7][9] , 
        \out_first_stage[7][8] , \out_first_stage[7][7] , 
        \out_first_stage[7][6] , \out_first_stage[7][5] , 
        \out_first_stage[7][4] , \out_first_stage[7][3] , 
        \out_first_stage[7][2] , \out_first_stage[7][1] , 
        \out_first_stage[7][0] }), .IN7({\out_first_stage[8][35] , 
        \out_first_stage[8][34] , \out_first_stage[8][33] , 
        \out_first_stage[8][32] , \out_first_stage[8][31] , 
        \out_first_stage[8][30] , \out_first_stage[8][29] , 
        \out_first_stage[8][28] , \out_first_stage[8][27] , 
        \out_first_stage[8][26] , \out_first_stage[8][25] , 
        \out_first_stage[8][24] , \out_first_stage[8][23] , 
        \out_first_stage[8][22] , \out_first_stage[8][21] , 
        \out_first_stage[8][20] , \out_first_stage[8][19] , 
        \out_first_stage[8][18] , \out_first_stage[8][17] , 
        \out_first_stage[8][16] , \out_first_stage[8][15] , 
        \out_first_stage[8][14] , \out_first_stage[8][13] , 
        \out_first_stage[8][12] , \out_first_stage[8][11] , 
        \out_first_stage[8][10] , \out_first_stage[8][9] , 
        \out_first_stage[8][8] , \out_first_stage[8][7] , 
        \out_first_stage[8][6] , \out_first_stage[8][5] , 
        \out_first_stage[8][4] , \out_first_stage[8][3] , 
        \out_first_stage[8][2] , \out_first_stage[8][1] , 
        \out_first_stage[8][0] }), .SEL(shift_pos[4:2]), .Y(out_second_stage)
         );
  MUX_8to1_N32_1 mux_third_stage ( .IN0({out_second_stage[35:14], 1'b0, 1'b0, 
        1'b0, 1'b0, out_second_stage[9:4]}), .IN1({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .IN2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .IN3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN4({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        out_second_stage[10], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, out_second_stage[0]}), .IN5({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, out_second_stage[11], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, out_second_stage[1]}), .IN6({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, out_second_stage[12], 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, out_second_stage[2]}), .IN7(
        {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        out_second_stage[13], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, out_second_stage[3]}), .SEL({n310, shift_pos[1:0]}), .Y(
        out_barrel) );
  MUX_2to1_N32_1 mux_out ( .IN0(out_control), .IN1(out_barrel), .SEL(n9), .Y(
        OUTPUT) );
  DLL_X1 \shift_pos_reg[4]  ( .D(B[4]), .GN(N0), .Q(shift_pos[4]) );
  DLL_X1 \shift_pos_reg[3]  ( .D(B[3]), .GN(N0), .Q(shift_pos[3]) );
  DLL_X1 \shift_pos_reg[2]  ( .D(B[2]), .GN(N0), .Q(shift_pos[2]) );
  DLL_X1 \shift_pos_reg[1]  ( .D(B[1]), .GN(N0), .Q(shift_pos[1]) );
  DLL_X1 \shift_pos_reg[0]  ( .D(B[0]), .GN(N0), .Q(shift_pos[0]) );
  DLH_X1 \out_control_reg[31]  ( .G(N0), .D(N1), .Q(out_control[31]) );
  DLH_X1 \out_control_reg[30]  ( .G(N0), .D(N1), .Q(out_control[30]) );
  DLH_X1 \out_control_reg[29]  ( .G(N0), .D(N1), .Q(out_control[29]) );
  DLH_X1 \out_control_reg[28]  ( .G(N0), .D(N1), .Q(out_control[28]) );
  DLH_X1 \out_control_reg[27]  ( .G(N0), .D(N1), .Q(out_control[27]) );
  DLH_X1 \out_control_reg[26]  ( .G(N0), .D(N1), .Q(out_control[26]) );
  DLH_X1 \out_control_reg[25]  ( .G(N0), .D(N1), .Q(out_control[25]) );
  DLH_X1 \out_control_reg[24]  ( .G(N0), .D(N1), .Q(out_control[24]) );
  DLH_X1 \out_control_reg[23]  ( .G(N0), .D(N1), .Q(out_control[23]) );
  DLH_X1 \out_control_reg[22]  ( .G(N0), .D(N1), .Q(out_control[22]) );
  DLH_X1 \out_control_reg[21]  ( .G(N0), .D(N1), .Q(out_control[21]) );
  DLH_X1 \out_control_reg[20]  ( .G(N0), .D(N1), .Q(out_control[20]) );
  DLH_X1 \out_control_reg[19]  ( .G(N0), .D(N1), .Q(out_control[19]) );
  DLH_X1 \out_control_reg[18]  ( .G(N0), .D(N1), .Q(out_control[18]) );
  DLH_X1 \out_control_reg[17]  ( .G(N0), .D(N1), .Q(out_control[17]) );
  DLH_X1 \out_control_reg[16]  ( .G(N0), .D(N1), .Q(out_control[16]) );
  DLH_X1 \out_control_reg[15]  ( .G(N0), .D(N1), .Q(out_control[15]) );
  DLH_X1 \out_control_reg[14]  ( .G(N0), .D(N1), .Q(out_control[14]) );
  DLH_X1 \out_control_reg[13]  ( .G(N0), .D(N1), .Q(out_control[13]) );
  DLH_X1 \out_control_reg[12]  ( .G(N0), .D(N1), .Q(out_control[12]) );
  DLH_X1 \out_control_reg[11]  ( .G(N0), .D(N1), .Q(out_control[11]) );
  DLH_X1 \out_control_reg[10]  ( .G(N0), .D(N1), .Q(out_control[10]) );
  DLH_X1 \out_control_reg[9]  ( .G(N0), .D(N1), .Q(out_control[9]) );
  DLH_X1 \out_control_reg[8]  ( .G(N0), .D(N1), .Q(out_control[8]) );
  DLH_X1 \out_control_reg[7]  ( .G(N0), .D(N1), .Q(out_control[7]) );
  DLH_X1 \out_control_reg[6]  ( .G(N0), .D(N1), .Q(out_control[6]) );
  DLH_X1 \out_control_reg[5]  ( .G(N0), .D(N1), .Q(out_control[5]) );
  DLH_X1 \out_control_reg[4]  ( .G(N0), .D(N1), .Q(out_control[4]) );
  DLH_X1 \out_control_reg[3]  ( .G(N0), .D(N1), .Q(out_control[3]) );
  DLH_X1 \out_control_reg[2]  ( .G(N0), .D(N1), .Q(out_control[2]) );
  DLH_X1 \out_control_reg[1]  ( .G(N0), .D(N1), .Q(out_control[1]) );
  DLH_X1 \out_control_reg[0]  ( .G(N0), .D(N1), .Q(out_control[0]) );
  AND2_X1 U3 ( .A1(n310), .A2(LOGIC_ARITH), .ZN(N1) );
  AND2_X2 U4 ( .A1(n319), .A2(n318), .ZN(n9) );
  NAND2_X2 U5 ( .A1(n9), .A2(n320), .ZN(N0) );
  BUF_X4 U6 ( .A(LOGIC_ARITH), .Z(n311) );
  BUF_X8 U7 ( .A(LEFT_RIGHT), .Z(n310) );
  NOR4_X1 U308 ( .A1(B[12]), .A2(B[6]), .A3(B[7]), .A4(B[15]), .ZN(n319) );
  OR4_X1 U309 ( .A1(B[9]), .A2(B[11]), .A3(B[8]), .A4(B[19]), .ZN(n317) );
  NOR4_X1 U310 ( .A1(B[13]), .A2(B[17]), .A3(B[28]), .A4(B[16]), .ZN(n315) );
  NOR4_X1 U311 ( .A1(B[22]), .A2(B[20]), .A3(B[21]), .A4(B[18]), .ZN(n314) );
  NOR4_X1 U312 ( .A1(B[25]), .A2(B[30]), .A3(B[23]), .A4(B[26]), .ZN(n313) );
  NOR4_X1 U313 ( .A1(B[27]), .A2(B[29]), .A3(B[31]), .A4(B[24]), .ZN(n312) );
  NAND4_X1 U314 ( .A1(n315), .A2(n314), .A3(n313), .A4(n312), .ZN(n316) );
  NOR4_X1 U315 ( .A1(B[10]), .A2(B[14]), .A3(n317), .A4(n316), .ZN(n318) );
  INV_X1 U316 ( .A(B[5]), .ZN(n320) );
endmodule


module PG_NETWORK_992 ( op1, op2, g, p );
  input op1, op2;
  output g, p;
  wire   n1;

  XNOR2_X1 U1 ( .A(op2), .B(n1), .ZN(p) );
  INV_X1 U2 ( .A(op1), .ZN(n1) );
  AND2_X1 U3 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_991 ( op1, op2, g, p );
  input op1, op2;
  output g, p;
  wire   n2;

  XNOR2_X1 U1 ( .A(op2), .B(n2), .ZN(p) );
  INV_X1 U2 ( .A(op1), .ZN(n2) );
  AND2_X1 U3 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_990 ( op1, op2, g, p );
  input op1, op2;
  output g, p;
  wire   n2;

  XNOR2_X1 U1 ( .A(op2), .B(n2), .ZN(p) );
  INV_X1 U2 ( .A(op1), .ZN(n2) );
  AND2_X1 U3 ( .A1(op1), .A2(op2), .ZN(g) );
endmodule


module PG_NETWORK_989 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  XOR2_X1 U1 ( .A(op1), .B(op2), .Z(p) );
  AND2_X1 U2 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_988 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_987 ( op1, op2, g, p );
  input op1, op2;
  output g, p;
  wire   n1;

  XNOR2_X1 U1 ( .A(op2), .B(n1), .ZN(p) );
  INV_X1 U2 ( .A(op1), .ZN(n1) );
  AND2_X1 U3 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_986 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_985 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  XOR2_X1 U1 ( .A(op1), .B(op2), .Z(p) );
  AND2_X1 U2 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_984 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_983 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_982 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_981 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_980 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_979 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_978 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_977 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  XOR2_X1 U1 ( .A(op1), .B(op2), .Z(p) );
  AND2_X1 U2 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_976 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_975 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_974 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_973 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_972 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_971 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_970 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_969 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_968 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_967 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_966 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_965 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_964 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_963 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_962 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_961 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module G_BLOCK_264 ( P_ik, G_ik, G_k1j, G_ij );
  input P_ik, G_ik, G_k1j;
  output G_ij;
  wire   n1, n2;

  INV_X1 U1 ( .A(G_ik), .ZN(n1) );
  NAND2_X1 U2 ( .A1(G_k1j), .A2(P_ik), .ZN(n2) );
  NAND2_X1 U3 ( .A1(n2), .A2(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_972 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij_BAR );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij_BAR;


  AND2_X1 U1 ( .A1(P_k1j), .A2(P_ik), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(G_k1j), .A(G_ik), .ZN(G_ij_BAR) );
endmodule


module PG_BLOCK_971 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_970 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_k1j), .A2(P_ik), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_969 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_968 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(G_k1j), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_967 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_966 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_965 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_964 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_963 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_962 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(G_k1j), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_961 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_960 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_959 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_958 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module G_BLOCK_263 ( P_ik, G_k1j, G_ij, G_ik_BAR );
  input P_ik, G_k1j, G_ik_BAR;
  output G_ij;
  wire   G_ik, n1;
  assign G_ik = G_ik_BAR;

  NAND2_X2 U1 ( .A1(n1), .A2(G_ik), .ZN(G_ij) );
  NAND2_X1 U2 ( .A1(G_k1j), .A2(P_ik), .ZN(n1) );
endmodule


module PG_BLOCK_957 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij_BAR );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij_BAR;


  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(G_ij_BAR) );
endmodule


module PG_BLOCK_956 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_955 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_954 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_953 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_952 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_951 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module G_BLOCK_262 ( P_ik, G_k1j, G_ij, G_ik_BAR );
  input P_ik, G_k1j, G_ik_BAR;
  output G_ij;
  wire   G_ik, n1;
  assign G_ik = G_ik_BAR;

  NAND2_X1 U1 ( .A1(n1), .A2(G_ik), .ZN(G_ij) );
  NAND2_X1 U2 ( .A1(G_k1j), .A2(P_ik), .ZN(n1) );
endmodule


module PG_BLOCK_950 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij_BAR );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij_BAR;


  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(G_ij_BAR) );
endmodule


module PG_BLOCK_949 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_948 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module G_BLOCK_261 ( P_ik, G_ik, G_k1j, G_ij );
  input P_ik, G_ik, G_k1j;
  output G_ij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(G_ij) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(G_k1j), .A(G_ik), .ZN(n1) );
endmodule


module G_BLOCK_260 ( P_ik, G_k1j, G_ij, G_ik_BAR );
  input P_ik, G_k1j, G_ik_BAR;
  output G_ij;
  wire   G_ik, n1;
  assign G_ik = G_ik_BAR;

  NAND2_X2 U1 ( .A1(n1), .A2(G_ik), .ZN(G_ij) );
  NAND2_X1 U2 ( .A1(G_k1j), .A2(P_ik), .ZN(n1) );
endmodule


module PG_BLOCK_947 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_946 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module G_BLOCK_259 ( P_ik, G_ik, G_k1j, G_ij );
  input P_ik, G_ik, G_k1j;
  output G_ij;
  wire   n1, n2;

  NAND2_X1 U1 ( .A1(n2), .A2(n1), .ZN(G_ij) );
  INV_X1 U2 ( .A(G_ik), .ZN(n1) );
  NAND2_X1 U3 ( .A1(G_k1j), .A2(P_ik), .ZN(n2) );
endmodule


module G_BLOCK_258 ( P_ik, G_ik, G_k1j, G_ij );
  input P_ik, G_ik, G_k1j;
  output G_ij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(G_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
endmodule


module G_BLOCK_257 ( P_ik, G_ik, G_k1j, G_ij );
  input P_ik, G_ik, G_k1j;
  output G_ij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(G_ij) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(G_k1j), .A(G_ik), .ZN(n1) );
endmodule


module G_BLOCK_256 ( P_ik, G_ik, G_k1j, G_ij );
  input P_ik, G_ik, G_k1j;
  output G_ij;
  wire   n1;

  AOI21_X1 U1 ( .B1(P_ik), .B2(G_k1j), .A(G_ik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(G_ij) );
endmodule


module CARRY_GENERATOR_Nbit32_1 ( A, B, Cin, Cout );
  input [31:0] A;
  input [31:0] B;
  output [8:0] Cout;
  input Cin;
  wire   Cin, n13, \p[4][3] , \p[4][2] , \p[3][3] , \p[3][2] , \p[3][1] ,
         \p[2][7] , \p[2][6] , \p[2][5] , \p[2][4] , \p[2][3] , \p[2][2] ,
         \p[2][1] , \p[1][15] , \p[1][14] , \p[1][13] , \p[1][12] , \p[1][11] ,
         \p[1][10] , \p[1][9] , \p[1][8] , \p[1][7] , \p[1][6] , \p[1][5] ,
         \p[1][4] , \p[1][3] , \p[1][2] , \p[1][1] , \p[0][32] , \p[0][31] ,
         \p[0][30] , \p[0][29] , \p[0][28] , \p[0][27] , \p[0][26] ,
         \p[0][25] , \p[0][24] , \p[0][23] , \p[0][22] , \p[0][21] ,
         \p[0][20] , \p[0][19] , \p[0][18] , \p[0][17] , \p[0][16] ,
         \p[0][15] , \p[0][14] , \p[0][13] , \p[0][12] , \p[0][11] ,
         \p[0][10] , \p[0][9] , \p[0][8] , \p[0][7] , \p[0][6] , \p[0][5] ,
         \p[0][4] , \p[0][3] , \p[0][2] , \p[0][1] , \g[4][3] , \g[4][2] ,
         \g[3][3] , \g[3][2] , \g[3][1] , \g[2][7] , \g[2][6] , \g[2][5] ,
         \g[2][4] , \g[2][3] , \g[2][2] , \g[2][1] , \g[1][15] , \g[1][14] ,
         \g[1][13] , \g[1][12] , \g[1][11] , \g[1][10] , \g[1][9] , \g[1][8] ,
         \g[1][7] , \g[1][6] , \g[1][5] , \g[1][4] , \g[1][3] , \g[1][2] ,
         \g[1][1] , \g[1][0] , \g[0][32] , \g[0][31] , \g[0][30] , \g[0][29] ,
         \g[0][28] , \g[0][27] , \g[0][26] , \g[0][25] , \g[0][24] ,
         \g[0][23] , \g[0][22] , \g[0][21] , \g[0][20] , \g[0][19] ,
         \g[0][18] , \g[0][17] , \g[0][16] , \g[0][15] , \g[0][14] ,
         \g[0][13] , \g[0][12] , \g[0][11] , \g[0][10] , \g[0][9] , \g[0][8] ,
         \g[0][7] , \g[0][6] , \g[0][5] , \g[0][4] , \g[0][3] , \g[0][2] ,
         \g[0][1] , n2, n3, n12;
  assign Cout[0] = Cin;

  PG_NETWORK_992 Block_PG_NET_1 ( .op1(A[0]), .op2(B[0]), .g(\g[0][1] ), .p(
        \p[0][1] ) );
  PG_NETWORK_991 Block_PG_NET_2 ( .op1(A[1]), .op2(B[1]), .g(\g[0][2] ), .p(
        \p[0][2] ) );
  PG_NETWORK_990 Block_PG_NET_3 ( .op1(A[2]), .op2(B[2]), .g(\g[0][3] ), .p(
        \p[0][3] ) );
  PG_NETWORK_989 Block_PG_NET_4 ( .op1(A[3]), .op2(B[3]), .g(\g[0][4] ), .p(
        \p[0][4] ) );
  PG_NETWORK_988 Block_PG_NET_5 ( .op1(A[4]), .op2(B[4]), .g(\g[0][5] ), .p(
        \p[0][5] ) );
  PG_NETWORK_987 Block_PG_NET_6 ( .op1(A[5]), .op2(B[5]), .g(\g[0][6] ), .p(
        \p[0][6] ) );
  PG_NETWORK_986 Block_PG_NET_7 ( .op1(A[6]), .op2(B[6]), .g(\g[0][7] ), .p(
        \p[0][7] ) );
  PG_NETWORK_985 Block_PG_NET_8 ( .op1(A[7]), .op2(B[7]), .g(\g[0][8] ), .p(
        \p[0][8] ) );
  PG_NETWORK_984 Block_PG_NET_9 ( .op1(A[8]), .op2(B[8]), .g(\g[0][9] ), .p(
        \p[0][9] ) );
  PG_NETWORK_983 Block_PG_NET_10 ( .op1(A[9]), .op2(B[9]), .g(\g[0][10] ), .p(
        \p[0][10] ) );
  PG_NETWORK_982 Block_PG_NET_11 ( .op1(A[10]), .op2(B[10]), .g(\g[0][11] ), 
        .p(\p[0][11] ) );
  PG_NETWORK_981 Block_PG_NET_12 ( .op1(A[11]), .op2(B[11]), .g(\g[0][12] ), 
        .p(\p[0][12] ) );
  PG_NETWORK_980 Block_PG_NET_13 ( .op1(A[12]), .op2(B[12]), .g(\g[0][13] ), 
        .p(\p[0][13] ) );
  PG_NETWORK_979 Block_PG_NET_14 ( .op1(A[13]), .op2(B[13]), .g(\g[0][14] ), 
        .p(\p[0][14] ) );
  PG_NETWORK_978 Block_PG_NET_15 ( .op1(A[14]), .op2(B[14]), .g(\g[0][15] ), 
        .p(\p[0][15] ) );
  PG_NETWORK_977 Block_PG_NET_16 ( .op1(A[15]), .op2(B[15]), .g(\g[0][16] ), 
        .p(\p[0][16] ) );
  PG_NETWORK_976 Block_PG_NET_17 ( .op1(A[16]), .op2(B[16]), .g(\g[0][17] ), 
        .p(\p[0][17] ) );
  PG_NETWORK_975 Block_PG_NET_18 ( .op1(A[17]), .op2(B[17]), .g(\g[0][18] ), 
        .p(\p[0][18] ) );
  PG_NETWORK_974 Block_PG_NET_19 ( .op1(A[18]), .op2(B[18]), .g(\g[0][19] ), 
        .p(\p[0][19] ) );
  PG_NETWORK_973 Block_PG_NET_20 ( .op1(A[19]), .op2(B[19]), .g(\g[0][20] ), 
        .p(\p[0][20] ) );
  PG_NETWORK_972 Block_PG_NET_21 ( .op1(A[20]), .op2(B[20]), .g(\g[0][21] ), 
        .p(\p[0][21] ) );
  PG_NETWORK_971 Block_PG_NET_22 ( .op1(A[21]), .op2(B[21]), .g(\g[0][22] ), 
        .p(\p[0][22] ) );
  PG_NETWORK_970 Block_PG_NET_23 ( .op1(A[22]), .op2(B[22]), .g(\g[0][23] ), 
        .p(\p[0][23] ) );
  PG_NETWORK_969 Block_PG_NET_24 ( .op1(A[23]), .op2(B[23]), .g(\g[0][24] ), 
        .p(\p[0][24] ) );
  PG_NETWORK_968 Block_PG_NET_25 ( .op1(A[24]), .op2(B[24]), .g(\g[0][25] ), 
        .p(\p[0][25] ) );
  PG_NETWORK_967 Block_PG_NET_26 ( .op1(A[25]), .op2(B[25]), .g(\g[0][26] ), 
        .p(\p[0][26] ) );
  PG_NETWORK_966 Block_PG_NET_27 ( .op1(A[26]), .op2(B[26]), .g(\g[0][27] ), 
        .p(\p[0][27] ) );
  PG_NETWORK_965 Block_PG_NET_28 ( .op1(A[27]), .op2(B[27]), .g(\g[0][28] ), 
        .p(\p[0][28] ) );
  PG_NETWORK_964 Block_PG_NET_29 ( .op1(A[28]), .op2(B[28]), .g(\g[0][29] ), 
        .p(\p[0][29] ) );
  PG_NETWORK_963 Block_PG_NET_30 ( .op1(A[29]), .op2(B[29]), .g(\g[0][30] ), 
        .p(\p[0][30] ) );
  PG_NETWORK_962 Block_PG_NET_31 ( .op1(A[30]), .op2(B[30]), .g(\g[0][31] ), 
        .p(\p[0][31] ) );
  PG_NETWORK_961 Block_PG_NET_32 ( .op1(A[31]), .op2(B[31]), .g(\g[0][32] ), 
        .p(\p[0][32] ) );
  G_BLOCK_264 g_1 ( .P_ik(\p[0][2] ), .G_ik(\g[0][2] ), .G_k1j(n12), .G_ij(
        \g[1][0] ) );
  PG_BLOCK_972 Block_Stage_ONE_1 ( .P_ik(\p[0][4] ), .G_ik(\g[0][4] ), .P_k1j(
        \p[0][3] ), .G_k1j(\g[0][3] ), .P_ij(\p[1][1] ), .G_ij_BAR(\g[1][1] )
         );
  PG_BLOCK_971 Block_Stage_ONE_2 ( .P_ik(\p[0][6] ), .G_ik(\g[0][6] ), .P_k1j(
        \p[0][5] ), .G_k1j(\g[0][5] ), .P_ij(\p[1][2] ), .G_ij(\g[1][2] ) );
  PG_BLOCK_970 Block_Stage_ONE_3 ( .P_ik(\p[0][8] ), .G_ik(\g[0][8] ), .P_k1j(
        \p[0][7] ), .G_k1j(\g[0][7] ), .P_ij(\p[1][3] ), .G_ij(\g[1][3] ) );
  PG_BLOCK_969 Block_Stage_ONE_4 ( .P_ik(\p[0][10] ), .G_ik(\g[0][10] ), 
        .P_k1j(\p[0][9] ), .G_k1j(\g[0][9] ), .P_ij(\p[1][4] ), .G_ij(
        \g[1][4] ) );
  PG_BLOCK_968 Block_Stage_ONE_5 ( .P_ik(\p[0][12] ), .G_ik(\g[0][12] ), 
        .P_k1j(\p[0][11] ), .G_k1j(\g[0][11] ), .P_ij(\p[1][5] ), .G_ij(
        \g[1][5] ) );
  PG_BLOCK_967 Block_Stage_ONE_6 ( .P_ik(\p[0][14] ), .G_ik(\g[0][14] ), 
        .P_k1j(\p[0][13] ), .G_k1j(\g[0][13] ), .P_ij(\p[1][6] ), .G_ij(
        \g[1][6] ) );
  PG_BLOCK_966 Block_Stage_ONE_7 ( .P_ik(\p[0][16] ), .G_ik(\g[0][16] ), 
        .P_k1j(\p[0][15] ), .G_k1j(\g[0][15] ), .P_ij(\p[1][7] ), .G_ij(
        \g[1][7] ) );
  PG_BLOCK_965 Block_Stage_ONE_8 ( .P_ik(\p[0][18] ), .G_ik(\g[0][18] ), 
        .P_k1j(\p[0][17] ), .G_k1j(\g[0][17] ), .P_ij(\p[1][8] ), .G_ij(
        \g[1][8] ) );
  PG_BLOCK_964 Block_Stage_ONE_9 ( .P_ik(\p[0][20] ), .G_ik(\g[0][20] ), 
        .P_k1j(\p[0][19] ), .G_k1j(\g[0][19] ), .P_ij(\p[1][9] ), .G_ij(
        \g[1][9] ) );
  PG_BLOCK_963 Block_Stage_ONE_10 ( .P_ik(\p[0][22] ), .G_ik(\g[0][22] ), 
        .P_k1j(\p[0][21] ), .G_k1j(\g[0][21] ), .P_ij(\p[1][10] ), .G_ij(
        \g[1][10] ) );
  PG_BLOCK_962 Block_Stage_ONE_11 ( .P_ik(\p[0][24] ), .G_ik(\g[0][24] ), 
        .P_k1j(\p[0][23] ), .G_k1j(\g[0][23] ), .P_ij(\p[1][11] ), .G_ij(
        \g[1][11] ) );
  PG_BLOCK_961 Block_Stage_ONE_12 ( .P_ik(\p[0][26] ), .G_ik(\g[0][26] ), 
        .P_k1j(\p[0][25] ), .G_k1j(\g[0][25] ), .P_ij(\p[1][12] ), .G_ij(
        \g[1][12] ) );
  PG_BLOCK_960 Block_Stage_ONE_13 ( .P_ik(\p[0][28] ), .G_ik(\g[0][28] ), 
        .P_k1j(\p[0][27] ), .G_k1j(\g[0][27] ), .P_ij(\p[1][13] ), .G_ij(
        \g[1][13] ) );
  PG_BLOCK_959 Block_Stage_ONE_14 ( .P_ik(\p[0][30] ), .G_ik(\g[0][30] ), 
        .P_k1j(\p[0][29] ), .G_k1j(\g[0][29] ), .P_ij(\p[1][14] ), .G_ij(
        \g[1][14] ) );
  PG_BLOCK_958 Block_Stage_ONE_15 ( .P_ik(\p[0][32] ), .G_ik(\g[0][32] ), 
        .P_k1j(\p[0][31] ), .G_k1j(\g[0][31] ), .P_ij(\p[1][15] ), .G_ij(
        \g[1][15] ) );
  G_BLOCK_263 g_2 ( .P_ik(\p[1][1] ), .G_k1j(\g[1][0] ), .G_ij(Cout[1]), 
        .G_ik_BAR(\g[1][1] ) );
  PG_BLOCK_957 Block_Stage_TWO_1 ( .P_ik(\p[1][3] ), .G_ik(\g[1][3] ), .P_k1j(
        \p[1][2] ), .G_k1j(\g[1][2] ), .P_ij(\p[2][1] ), .G_ij_BAR(\g[2][1] )
         );
  PG_BLOCK_956 Block_Stage_TWO_2 ( .P_ik(\p[1][5] ), .G_ik(\g[1][5] ), .P_k1j(
        \p[1][4] ), .G_k1j(\g[1][4] ), .P_ij(\p[2][2] ), .G_ij(\g[2][2] ) );
  PG_BLOCK_955 Block_Stage_TWO_3 ( .P_ik(\p[1][7] ), .G_ik(\g[1][7] ), .P_k1j(
        \p[1][6] ), .G_k1j(\g[1][6] ), .P_ij(\p[2][3] ), .G_ij(\g[2][3] ) );
  PG_BLOCK_954 Block_Stage_TWO_4 ( .P_ik(\p[1][9] ), .G_ik(\g[1][9] ), .P_k1j(
        \p[1][8] ), .G_k1j(\g[1][8] ), .P_ij(\p[2][4] ), .G_ij(\g[2][4] ) );
  PG_BLOCK_953 Block_Stage_TWO_5 ( .P_ik(\p[1][11] ), .G_ik(\g[1][11] ), 
        .P_k1j(\p[1][10] ), .G_k1j(\g[1][10] ), .P_ij(\p[2][5] ), .G_ij(
        \g[2][5] ) );
  PG_BLOCK_952 Block_Stage_TWO_6 ( .P_ik(\p[1][13] ), .G_ik(\g[1][13] ), 
        .P_k1j(\p[1][12] ), .G_k1j(\g[1][12] ), .P_ij(\p[2][6] ), .G_ij(
        \g[2][6] ) );
  PG_BLOCK_951 Block_Stage_TWO_7 ( .P_ik(\p[1][15] ), .G_ik(\g[1][15] ), 
        .P_k1j(\p[1][14] ), .G_k1j(\g[1][14] ), .P_ij(\p[2][7] ), .G_ij(
        \g[2][7] ) );
  G_BLOCK_262 g_3 ( .P_ik(\p[2][1] ), .G_k1j(Cout[1]), .G_ij(n13), .G_ik_BAR(
        \g[2][1] ) );
  PG_BLOCK_950 Block_Stage_THREE_1 ( .P_ik(\p[2][3] ), .G_ik(\g[2][3] ), 
        .P_k1j(\p[2][2] ), .G_k1j(\g[2][2] ), .P_ij(\p[3][1] ), .G_ij_BAR(
        \g[3][1] ) );
  PG_BLOCK_949 Block_Stage_THREE_2 ( .P_ik(\p[2][5] ), .G_ik(\g[2][5] ), 
        .P_k1j(\p[2][4] ), .G_k1j(\g[2][4] ), .P_ij(\p[3][2] ), .G_ij(
        \g[3][2] ) );
  PG_BLOCK_948 Block_Stage_THREE_3 ( .P_ik(\p[2][7] ), .G_ik(\g[2][7] ), 
        .P_k1j(\p[2][6] ), .G_k1j(\g[2][6] ), .P_ij(\p[3][3] ), .G_ij(
        \g[3][3] ) );
  G_BLOCK_261 g_4_c12_c16_0 ( .P_ik(\p[2][2] ), .G_ik(\g[2][2] ), .G_k1j(n3), 
        .G_ij(Cout[3]) );
  G_BLOCK_260 g_4_c12_c16_1 ( .P_ik(\p[3][1] ), .G_k1j(n13), .G_ij(Cout[4]), 
        .G_ik_BAR(\g[3][1] ) );
  PG_BLOCK_947 Block_stage_FOUR_2_0 ( .P_ik(\p[2][6] ), .G_ik(\g[2][6] ), 
        .P_k1j(\p[3][2] ), .G_k1j(\g[3][2] ), .P_ij(\p[4][2] ), .G_ij(
        \g[4][2] ) );
  PG_BLOCK_946 Block_stage_FOUR_2_1 ( .P_ik(\p[3][3] ), .G_ik(\g[3][3] ), 
        .P_k1j(\p[3][2] ), .G_k1j(\g[3][2] ), .P_ij(\p[4][3] ), .G_ij(
        \g[4][3] ) );
  G_BLOCK_259 Block_stage_FIVE_4 ( .P_ik(\p[2][4] ), .G_ik(\g[2][4] ), .G_k1j(
        Cout[4]), .G_ij(Cout[5]) );
  G_BLOCK_258 Block_stage_FIVE_5 ( .P_ik(\p[3][2] ), .G_ik(\g[3][2] ), .G_k1j(
        Cout[4]), .G_ij(Cout[6]) );
  G_BLOCK_257 Block_stage_FIVE_6 ( .P_ik(\p[4][2] ), .G_ik(\g[4][2] ), .G_k1j(
        Cout[4]), .G_ij(Cout[7]) );
  G_BLOCK_256 Block_stage_FIVE_7 ( .P_ik(\p[4][3] ), .G_ik(\g[4][3] ), .G_k1j(
        Cout[4]), .G_ij(Cout[8]) );
  AOI21_X1 U1 ( .B1(\p[0][1] ), .B2(Cin), .A(\g[0][1] ), .ZN(n2) );
  INV_X1 U2 ( .A(n2), .ZN(n12) );
  BUF_X1 U3 ( .A(n13), .Z(n3) );
  BUF_X2 U4 ( .A(n13), .Z(Cout[2]) );
endmodule


module FA_1984 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1983 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1982 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(Ci), .CI(B), .CO(Co), .S(S) );
endmodule


module FA_1981 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_496 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1984 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1983 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1982 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1981 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1980 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_1979 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1978 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1977 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_495 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1980 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1979 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1978 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1977 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_248 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U3 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U4 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
endmodule


module carry_select_block_N4_248 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_496 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_495 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_248 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_1976 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1975 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(Ci), .CI(B), .CO(Co), .S(S) );
endmodule


module FA_1974 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1973 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_494 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1976 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1975 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1974 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1973 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1972 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_1971 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1970 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1969 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_493 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1972 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1971 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1970 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1969 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_247 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U3 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U4 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
endmodule


module carry_select_block_N4_247 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_494 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_493 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_247 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_1968 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1967 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1966 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1965 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_492 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1968 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1967 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1966 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1965 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1964 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_1963 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1962 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1961 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_491 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1964 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1963 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1962 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1961 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_246 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U3 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U4 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
endmodule


module carry_select_block_N4_246 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_492 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_491 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_246 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_1960 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1959 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1958 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1957 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_490 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1960 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1959 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1958 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1957 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1956 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_1955 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1954 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1953 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_489 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1956 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1955 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1954 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1953 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_245 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U3 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U4 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
endmodule


module carry_select_block_N4_245 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_490 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_489 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_245 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_1952 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1951 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1950 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1949 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n2) );
  XNOR2_X1 U2 ( .A(n2), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_488 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1952 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1951 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1950 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1949 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1948 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_1947 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1946 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1945 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n2) );
  XNOR2_X1 U2 ( .A(n2), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_487 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1948 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1947 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1946 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1945 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_244 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U3 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U4 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
endmodule


module carry_select_block_N4_244 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_488 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_487 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_244 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_1944 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1943 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1942 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1941 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_486 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1944 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1943 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1942 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1941 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1940 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_1939 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1938 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1937 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_485 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1940 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1939 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1938 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1937 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_243 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;
  wire   n1, n2;

  INV_X1 U1 ( .A(IN0[3]), .ZN(n2) );
  NAND2_X1 U2 ( .A1(SEL), .A2(IN1[3]), .ZN(n1) );
  OAI21_X1 U3 ( .B1(SEL), .B2(n2), .A(n1), .ZN(Y[3]) );
  MUX2_X1 U4 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U5 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U6 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
endmodule


module carry_select_block_N4_243 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_486 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_485 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_243 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_1936 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1935 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1934 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1933 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_484 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1936 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1935 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1934 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1933 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1932 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_1931 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1930 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1929 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_483 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1932 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1931 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1930 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1929 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_242 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U3 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U4 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
endmodule


module carry_select_block_N4_242 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_484 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_483 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_242 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_1928 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1927 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1926 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1925 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_482 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1928 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1927 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1926 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1925 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1924 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_1923 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1922 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1921 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_481 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1924 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1923 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1922 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1921 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_241 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U3 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U4 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
endmodule


module carry_select_block_N4_241 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_482 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_481 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_241 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module SUMGENERATOR_Nblocks8_bits_per_block4_1 ( A, B, CARRY_SELECT, SUM );
  input [31:0] A;
  input [31:0] B;
  input [7:0] CARRY_SELECT;
  output [31:0] SUM;


  carry_select_block_N4_248 block_n_1 ( .A(A[3:0]), .B(B[3:0]), .S(SUM[3:0]), 
        .Ci(CARRY_SELECT[0]) );
  carry_select_block_N4_247 block_n_2 ( .A(A[7:4]), .B(B[7:4]), .S(SUM[7:4]), 
        .Ci(CARRY_SELECT[1]) );
  carry_select_block_N4_246 block_n_3 ( .A(A[11:8]), .B(B[11:8]), .S(SUM[11:8]), .Ci(CARRY_SELECT[2]) );
  carry_select_block_N4_245 block_n_4 ( .A(A[15:12]), .B(B[15:12]), .S(
        SUM[15:12]), .Ci(CARRY_SELECT[3]) );
  carry_select_block_N4_244 block_n_5 ( .A(A[19:16]), .B(B[19:16]), .S(
        SUM[19:16]), .Ci(CARRY_SELECT[4]) );
  carry_select_block_N4_243 block_n_6 ( .A(A[23:20]), .B(B[23:20]), .S(
        SUM[23:20]), .Ci(CARRY_SELECT[5]) );
  carry_select_block_N4_242 block_n_7 ( .A(A[27:24]), .B(B[27:24]), .S(
        SUM[27:24]), .Ci(CARRY_SELECT[6]) );
  carry_select_block_N4_241 block_n_8 ( .A(A[31:28]), .B(B[31:28]), .S(
        SUM[31:28]), .Ci(CARRY_SELECT[7]) );
endmodule


module ADDER_P4_N_BIT32_1 ( A, B, add_sub, Cout, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input add_sub;
  output Cout;
  wire   n1, n2, n11, n12, n13, n14, n15;
  wire   [31:0] B_xor;
  wire   [7:0] tmp_co;

  CARRY_GENERATOR_Nbit32_1 CLA_SPARSE_TREE ( .A(A), .B(B_xor), .Cin(n11), 
        .Cout({Cout, tmp_co}) );
  SUMGENERATOR_Nblocks8_bits_per_block4_1 CSA ( .A(A), .B({B_xor[31:4], n2, 
        B_xor[2], n13, B_xor[0]}), .CARRY_SELECT(tmp_co), .SUM(SUM) );
  XOR2_X1 U1 ( .A(B[3]), .B(n12), .Z(B_xor[3]) );
  XOR2_X1 U2 ( .A(B[2]), .B(n12), .Z(B_xor[2]) );
  INV_X1 U3 ( .A(n15), .ZN(n1) );
  XOR2_X1 U4 ( .A(B[5]), .B(n12), .Z(B_xor[5]) );
  BUF_X1 U5 ( .A(B_xor[3]), .Z(n2) );
  BUF_X2 U6 ( .A(add_sub), .Z(n12) );
  XNOR2_X2 U7 ( .A(B[0]), .B(n15), .ZN(B_xor[0]) );
  INV_X1 U8 ( .A(n15), .ZN(n11) );
  XNOR2_X1 U9 ( .A(n1), .B(n14), .ZN(n13) );
  XOR2_X1 U10 ( .A(n12), .B(B[9]), .Z(B_xor[9]) );
  XOR2_X1 U11 ( .A(n12), .B(B[11]), .Z(B_xor[11]) );
  XOR2_X1 U12 ( .A(n1), .B(B[12]), .Z(B_xor[12]) );
  XOR2_X1 U13 ( .A(n12), .B(B[13]), .Z(B_xor[13]) );
  XOR2_X1 U14 ( .A(n12), .B(B[14]), .Z(B_xor[14]) );
  XOR2_X1 U15 ( .A(n12), .B(B[15]), .Z(B_xor[15]) );
  XOR2_X1 U16 ( .A(n12), .B(B[6]), .Z(B_xor[6]) );
  XOR2_X1 U17 ( .A(n12), .B(B[7]), .Z(B_xor[7]) );
  INV_X1 U18 ( .A(add_sub), .ZN(n15) );
  XNOR2_X1 U19 ( .A(n1), .B(n14), .ZN(B_xor[1]) );
  INV_X1 U20 ( .A(B[1]), .ZN(n14) );
  XOR2_X1 U21 ( .A(n12), .B(B[10]), .Z(B_xor[10]) );
  XOR2_X1 U22 ( .A(n1), .B(B[16]), .Z(B_xor[16]) );
  XOR2_X1 U23 ( .A(n1), .B(B[17]), .Z(B_xor[17]) );
  XOR2_X1 U24 ( .A(tmp_co[0]), .B(B[18]), .Z(B_xor[18]) );
  XOR2_X1 U25 ( .A(n12), .B(B[19]), .Z(B_xor[19]) );
  XOR2_X1 U26 ( .A(tmp_co[0]), .B(B[20]), .Z(B_xor[20]) );
  XOR2_X1 U27 ( .A(n12), .B(B[21]), .Z(B_xor[21]) );
  XOR2_X1 U28 ( .A(n1), .B(B[22]), .Z(B_xor[22]) );
  XOR2_X1 U29 ( .A(n12), .B(B[23]), .Z(B_xor[23]) );
  XOR2_X1 U30 ( .A(n11), .B(B[24]), .Z(B_xor[24]) );
  XOR2_X1 U31 ( .A(n1), .B(B[25]), .Z(B_xor[25]) );
  XOR2_X1 U32 ( .A(n11), .B(B[26]), .Z(B_xor[26]) );
  XOR2_X1 U33 ( .A(n1), .B(B[27]), .Z(B_xor[27]) );
  XOR2_X1 U34 ( .A(n11), .B(B[28]), .Z(B_xor[28]) );
  XOR2_X1 U35 ( .A(n11), .B(B[29]), .Z(B_xor[29]) );
  XOR2_X1 U36 ( .A(n11), .B(B[30]), .Z(B_xor[30]) );
  XOR2_X1 U37 ( .A(n11), .B(B[31]), .Z(B_xor[31]) );
  XOR2_X1 U38 ( .A(n12), .B(B[4]), .Z(B_xor[4]) );
  XOR2_X1 U39 ( .A(n1), .B(B[8]), .Z(B_xor[8]) );
endmodule


module LOGIC_BLOCK_N32 ( SUM, C_OUT, A, B, A_GEU_B, A_GE_B, A_GT_B, A_GTU_B, 
        A_LEU_B, A_LE_B, A_LT_B, A_LTU_B, A_NE_B, A_EQ_B, NOT_A, A_AND_B, 
        A_XOR_B, A_OR_B );
  input [31:0] SUM;
  input [31:0] A;
  input [31:0] B;
  output [31:0] A_GEU_B;
  output [31:0] A_GE_B;
  output [31:0] A_GT_B;
  output [31:0] A_GTU_B;
  output [31:0] A_LEU_B;
  output [31:0] A_LE_B;
  output [31:0] A_LT_B;
  output [31:0] A_LTU_B;
  output [31:0] A_NE_B;
  output [31:0] A_EQ_B;
  output [31:0] NOT_A;
  output [31:0] A_AND_B;
  output [31:0] A_XOR_B;
  output [31:0] A_OR_B;
  input C_OUT;
  wire   C_OUT, n101, n1, n2, n3, n4, n5, n15, n16, n17, n18, n31, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100;
  assign A_GEU_B[0] = C_OUT;

  INV_X1 U2 ( .A(B[13]), .ZN(n1) );
  NAND2_X1 U3 ( .A1(NOT_A[13]), .A2(n1), .ZN(A_OR_B[13]) );
  INV_X1 U4 ( .A(A_OR_B[13]), .ZN(n2) );
  NOR2_X1 U5 ( .A1(NOT_A[13]), .A2(n1), .ZN(A_AND_B[13]) );
  NOR2_X1 U6 ( .A1(n2), .A2(A_AND_B[13]), .ZN(A_XOR_B[13]) );
  INV_X1 U7 ( .A(n93), .ZN(A_OR_B[30]) );
  NOR2_X1 U8 ( .A1(n93), .A2(A_AND_B[30]), .ZN(A_XOR_B[30]) );
  INV_X1 U9 ( .A(A[30]), .ZN(NOT_A[30]) );
  NAND2_X1 U10 ( .A1(n101), .A2(C_OUT), .ZN(n3) );
  AND4_X1 U11 ( .A1(n49), .A2(n51), .A3(n50), .A4(n64), .ZN(n5) );
  NAND2_X1 U12 ( .A1(n4), .A2(n5), .ZN(n101) );
  AND4_X1 U13 ( .A1(n65), .A2(n67), .A3(n52), .A4(n66), .ZN(n4) );
  XNOR2_X1 U14 ( .A(n3), .B(n70), .ZN(A_LE_B[0]) );
  NAND2_X1 U15 ( .A1(n101), .A2(C_OUT), .ZN(A_LEU_B[0]) );
  INV_X1 U16 ( .A(C_OUT), .ZN(n68) );
  AND2_X1 U17 ( .A1(B[31]), .A2(A[31]), .ZN(A_AND_B[31]) );
  AOI21_X1 U18 ( .B1(n68), .B2(n70), .A(n69), .ZN(A_GE_B[0]) );
  NOR2_X1 U19 ( .A1(n68), .A2(n70), .ZN(n69) );
  INV_X1 U20 ( .A(SUM[24]), .ZN(n64) );
  NOR2_X1 U21 ( .A1(SUM[28]), .A2(SUM[27]), .ZN(n51) );
  NOR2_X1 U22 ( .A1(SUM[30]), .A2(SUM[29]), .ZN(n52) );
  NAND2_X1 U23 ( .A1(n62), .A2(n61), .ZN(n63) );
  NOR2_X1 U24 ( .A1(SUM[13]), .A2(SUM[12]), .ZN(n61) );
  NOR2_X1 U25 ( .A1(SUM[19]), .A2(SUM[18]), .ZN(n62) );
  NOR3_X1 U26 ( .A1(n60), .A2(SUM[17]), .A3(SUM[16]), .ZN(n67) );
  NAND4_X1 U27 ( .A1(n17), .A2(n16), .A3(n59), .A4(n15), .ZN(n60) );
  AND2_X1 U28 ( .A1(n57), .A2(n58), .ZN(n15) );
  NOR2_X1 U29 ( .A1(SUM[10]), .A2(SUM[9]), .ZN(n58) );
  NOR3_X1 U30 ( .A1(SUM[8]), .A2(SUM[6]), .A3(SUM[2]), .ZN(n57) );
  NOR4_X1 U31 ( .A1(SUM[11]), .A2(n56), .A3(SUM[3]), .A4(SUM[7]), .ZN(n59) );
  NOR2_X1 U32 ( .A1(SUM[1]), .A2(SUM[0]), .ZN(n53) );
  INV_X1 U33 ( .A(SUM[5]), .ZN(n54) );
  INV_X1 U34 ( .A(SUM[4]), .ZN(n55) );
  INV_X1 U35 ( .A(SUM[15]), .ZN(n16) );
  INV_X1 U36 ( .A(SUM[14]), .ZN(n17) );
  NOR2_X1 U37 ( .A1(SUM[22]), .A2(SUM[21]), .ZN(n65) );
  INV_X1 U38 ( .A(A_XOR_B[31]), .ZN(n70) );
  OR2_X1 U39 ( .A1(B[31]), .A2(A[31]), .ZN(A_OR_B[31]) );
  AND2_X1 U40 ( .A1(n101), .A2(n68), .ZN(A_LTU_B[0]) );
  INV_X1 U41 ( .A(NOT_A[24]), .ZN(n18) );
  INV_X1 U42 ( .A(A[24]), .ZN(NOT_A[24]) );
  INV_X1 U43 ( .A(A[25]), .ZN(NOT_A[25]) );
  NOR2_X1 U44 ( .A1(SUM[26]), .A2(SUM[25]), .ZN(n50) );
  NOR2_X1 U45 ( .A1(SUM[31]), .A2(SUM[20]), .ZN(n49) );
  NOR2_X1 U46 ( .A1(n63), .A2(SUM[23]), .ZN(n66) );
  AND2_X1 U47 ( .A1(A_LE_B[0]), .A2(n101), .ZN(A_LT_B[0]) );
  INV_X1 U48 ( .A(n101), .ZN(A_EQ_B[0]) );
  AND2_X1 U49 ( .A1(n101), .A2(A_GE_B[0]), .ZN(A_GT_B[0]) );
  INV_X1 U50 ( .A(A[0]), .ZN(NOT_A[0]) );
  INV_X1 U51 ( .A(A[1]), .ZN(NOT_A[1]) );
  INV_X1 U52 ( .A(A[2]), .ZN(NOT_A[2]) );
  INV_X1 U53 ( .A(A[3]), .ZN(NOT_A[3]) );
  INV_X1 U54 ( .A(A[4]), .ZN(NOT_A[4]) );
  INV_X1 U55 ( .A(A[5]), .ZN(NOT_A[5]) );
  INV_X1 U56 ( .A(A[6]), .ZN(NOT_A[6]) );
  INV_X1 U57 ( .A(A[7]), .ZN(NOT_A[7]) );
  INV_X1 U58 ( .A(A[8]), .ZN(NOT_A[8]) );
  INV_X1 U59 ( .A(A[9]), .ZN(NOT_A[9]) );
  INV_X1 U60 ( .A(NOT_A[10]), .ZN(n31) );
  INV_X1 U61 ( .A(A[10]), .ZN(NOT_A[10]) );
  INV_X1 U62 ( .A(A[11]), .ZN(NOT_A[11]) );
  INV_X1 U63 ( .A(A[12]), .ZN(NOT_A[12]) );
  INV_X1 U64 ( .A(A[13]), .ZN(NOT_A[13]) );
  INV_X1 U65 ( .A(A[14]), .ZN(NOT_A[14]) );
  INV_X1 U66 ( .A(A[15]), .ZN(NOT_A[15]) );
  INV_X1 U67 ( .A(A[16]), .ZN(NOT_A[16]) );
  INV_X1 U68 ( .A(A[17]), .ZN(NOT_A[17]) );
  INV_X1 U69 ( .A(A[18]), .ZN(NOT_A[18]) );
  INV_X1 U70 ( .A(A[19]), .ZN(NOT_A[19]) );
  INV_X1 U71 ( .A(A[20]), .ZN(NOT_A[20]) );
  INV_X1 U72 ( .A(A[21]), .ZN(NOT_A[21]) );
  INV_X1 U73 ( .A(A[22]), .ZN(NOT_A[22]) );
  INV_X1 U74 ( .A(A[23]), .ZN(NOT_A[23]) );
  INV_X1 U75 ( .A(A[26]), .ZN(NOT_A[26]) );
  INV_X1 U76 ( .A(A[27]), .ZN(NOT_A[27]) );
  INV_X1 U77 ( .A(A[28]), .ZN(NOT_A[28]) );
  XOR2_X1 U78 ( .A(A[31]), .B(B[31]), .Z(A_XOR_B[31]) );
  NAND3_X1 U79 ( .A1(n55), .A2(n54), .A3(n53), .ZN(n56) );
  AND2_X1 U80 ( .A1(B[0]), .A2(A[0]), .ZN(A_AND_B[0]) );
  AND2_X1 U81 ( .A1(B[10]), .A2(n31), .ZN(A_AND_B[10]) );
  AND2_X1 U82 ( .A1(B[11]), .A2(A[11]), .ZN(A_AND_B[11]) );
  AND2_X1 U83 ( .A1(B[12]), .A2(A[12]), .ZN(A_AND_B[12]) );
  AND2_X1 U84 ( .A1(B[14]), .A2(A[14]), .ZN(A_AND_B[14]) );
  AND2_X1 U85 ( .A1(B[15]), .A2(A[15]), .ZN(A_AND_B[15]) );
  AND2_X1 U86 ( .A1(B[16]), .A2(A[16]), .ZN(A_AND_B[16]) );
  AND2_X1 U87 ( .A1(B[17]), .A2(A[17]), .ZN(A_AND_B[17]) );
  AND2_X1 U88 ( .A1(B[18]), .A2(A[18]), .ZN(A_AND_B[18]) );
  AND2_X1 U89 ( .A1(B[19]), .A2(A[19]), .ZN(A_AND_B[19]) );
  AND2_X1 U90 ( .A1(B[1]), .A2(A[1]), .ZN(A_AND_B[1]) );
  AND2_X1 U91 ( .A1(B[20]), .A2(A[20]), .ZN(A_AND_B[20]) );
  AND2_X1 U92 ( .A1(B[21]), .A2(A[21]), .ZN(A_AND_B[21]) );
  AND2_X1 U93 ( .A1(B[22]), .A2(A[22]), .ZN(A_AND_B[22]) );
  AND2_X1 U94 ( .A1(B[23]), .A2(A[23]), .ZN(A_AND_B[23]) );
  AND2_X1 U95 ( .A1(B[24]), .A2(n18), .ZN(A_AND_B[24]) );
  AND2_X1 U96 ( .A1(B[25]), .A2(A[25]), .ZN(A_AND_B[25]) );
  AND2_X1 U97 ( .A1(B[26]), .A2(A[26]), .ZN(A_AND_B[26]) );
  AND2_X1 U98 ( .A1(B[27]), .A2(A[27]), .ZN(A_AND_B[27]) );
  AND2_X1 U99 ( .A1(B[28]), .A2(A[28]), .ZN(A_AND_B[28]) );
  INV_X1 U100 ( .A(A[29]), .ZN(NOT_A[29]) );
  AND2_X1 U101 ( .A1(B[29]), .A2(A[29]), .ZN(A_AND_B[29]) );
  AND2_X1 U102 ( .A1(B[2]), .A2(A[2]), .ZN(A_AND_B[2]) );
  AND2_X1 U103 ( .A1(B[30]), .A2(A[30]), .ZN(A_AND_B[30]) );
  INV_X1 U104 ( .A(A[31]), .ZN(NOT_A[31]) );
  AND2_X1 U105 ( .A1(B[3]), .A2(A[3]), .ZN(A_AND_B[3]) );
  AND2_X1 U106 ( .A1(B[4]), .A2(A[4]), .ZN(A_AND_B[4]) );
  AND2_X1 U107 ( .A1(B[5]), .A2(A[5]), .ZN(A_AND_B[5]) );
  AND2_X1 U108 ( .A1(B[6]), .A2(A[6]), .ZN(A_AND_B[6]) );
  AND2_X1 U109 ( .A1(B[7]), .A2(A[7]), .ZN(A_AND_B[7]) );
  AND2_X1 U110 ( .A1(B[8]), .A2(A[8]), .ZN(A_AND_B[8]) );
  AND2_X1 U111 ( .A1(B[9]), .A2(A[9]), .ZN(A_AND_B[9]) );
  NOR2_X1 U112 ( .A1(B[0]), .A2(A[0]), .ZN(n71) );
  INV_X1 U113 ( .A(n71), .ZN(A_OR_B[0]) );
  NOR2_X1 U114 ( .A1(B[10]), .A2(n31), .ZN(n72) );
  INV_X1 U115 ( .A(n72), .ZN(A_OR_B[10]) );
  NOR2_X1 U116 ( .A1(B[11]), .A2(A[11]), .ZN(n73) );
  INV_X1 U117 ( .A(n73), .ZN(A_OR_B[11]) );
  NOR2_X1 U118 ( .A1(B[12]), .A2(A[12]), .ZN(n74) );
  INV_X1 U119 ( .A(n74), .ZN(A_OR_B[12]) );
  NOR2_X1 U120 ( .A1(B[14]), .A2(A[14]), .ZN(n75) );
  INV_X1 U121 ( .A(n75), .ZN(A_OR_B[14]) );
  NOR2_X1 U122 ( .A1(B[15]), .A2(A[15]), .ZN(n76) );
  INV_X1 U123 ( .A(n76), .ZN(A_OR_B[15]) );
  NOR2_X1 U124 ( .A1(B[16]), .A2(A[16]), .ZN(n77) );
  INV_X1 U125 ( .A(n77), .ZN(A_OR_B[16]) );
  NOR2_X1 U126 ( .A1(B[17]), .A2(A[17]), .ZN(n78) );
  INV_X1 U127 ( .A(n78), .ZN(A_OR_B[17]) );
  NOR2_X1 U128 ( .A1(B[18]), .A2(A[18]), .ZN(n79) );
  INV_X1 U129 ( .A(n79), .ZN(A_OR_B[18]) );
  NOR2_X1 U130 ( .A1(B[19]), .A2(A[19]), .ZN(n80) );
  INV_X1 U131 ( .A(n80), .ZN(A_OR_B[19]) );
  NOR2_X1 U132 ( .A1(B[1]), .A2(A[1]), .ZN(n81) );
  INV_X1 U133 ( .A(n81), .ZN(A_OR_B[1]) );
  NOR2_X1 U134 ( .A1(B[20]), .A2(A[20]), .ZN(n82) );
  INV_X1 U135 ( .A(n82), .ZN(A_OR_B[20]) );
  NOR2_X1 U136 ( .A1(B[21]), .A2(A[21]), .ZN(n83) );
  INV_X1 U137 ( .A(n83), .ZN(A_OR_B[21]) );
  NOR2_X1 U138 ( .A1(B[22]), .A2(A[22]), .ZN(n84) );
  INV_X1 U139 ( .A(n84), .ZN(A_OR_B[22]) );
  NOR2_X1 U140 ( .A1(B[23]), .A2(A[23]), .ZN(n85) );
  INV_X1 U141 ( .A(n85), .ZN(A_OR_B[23]) );
  NOR2_X1 U142 ( .A1(B[24]), .A2(n18), .ZN(n86) );
  INV_X1 U143 ( .A(n86), .ZN(A_OR_B[24]) );
  NOR2_X1 U144 ( .A1(B[25]), .A2(A[25]), .ZN(n87) );
  INV_X1 U145 ( .A(n87), .ZN(A_OR_B[25]) );
  NOR2_X1 U146 ( .A1(B[26]), .A2(A[26]), .ZN(n88) );
  INV_X1 U147 ( .A(n88), .ZN(A_OR_B[26]) );
  NOR2_X1 U148 ( .A1(B[27]), .A2(A[27]), .ZN(n89) );
  INV_X1 U149 ( .A(n89), .ZN(A_OR_B[27]) );
  NOR2_X1 U150 ( .A1(B[28]), .A2(A[28]), .ZN(n90) );
  INV_X1 U151 ( .A(n90), .ZN(A_OR_B[28]) );
  NOR2_X1 U152 ( .A1(B[29]), .A2(A[29]), .ZN(n91) );
  INV_X1 U153 ( .A(n91), .ZN(A_OR_B[29]) );
  NOR2_X1 U154 ( .A1(A[2]), .A2(B[2]), .ZN(n92) );
  INV_X1 U155 ( .A(n92), .ZN(A_OR_B[2]) );
  NOR2_X1 U156 ( .A1(B[30]), .A2(A[30]), .ZN(n93) );
  NOR2_X1 U157 ( .A1(A[3]), .A2(B[3]), .ZN(n94) );
  INV_X1 U158 ( .A(n94), .ZN(A_OR_B[3]) );
  NOR2_X1 U159 ( .A1(B[4]), .A2(A[4]), .ZN(n95) );
  INV_X1 U160 ( .A(n95), .ZN(A_OR_B[4]) );
  NOR2_X1 U161 ( .A1(B[5]), .A2(A[5]), .ZN(n96) );
  INV_X1 U162 ( .A(n96), .ZN(A_OR_B[5]) );
  NOR2_X1 U163 ( .A1(B[6]), .A2(A[6]), .ZN(n97) );
  INV_X1 U164 ( .A(n97), .ZN(A_OR_B[6]) );
  NOR2_X1 U165 ( .A1(B[7]), .A2(A[7]), .ZN(n98) );
  INV_X1 U166 ( .A(n98), .ZN(A_OR_B[7]) );
  NOR2_X1 U167 ( .A1(B[8]), .A2(A[8]), .ZN(n99) );
  INV_X1 U168 ( .A(n99), .ZN(A_OR_B[8]) );
  NOR2_X1 U169 ( .A1(B[9]), .A2(A[9]), .ZN(n100) );
  INV_X1 U170 ( .A(n100), .ZN(A_OR_B[9]) );
  NOR2_X1 U171 ( .A1(n71), .A2(A_AND_B[0]), .ZN(A_XOR_B[0]) );
  NOR2_X1 U172 ( .A1(n72), .A2(A_AND_B[10]), .ZN(A_XOR_B[10]) );
  NOR2_X1 U173 ( .A1(n73), .A2(A_AND_B[11]), .ZN(A_XOR_B[11]) );
  NOR2_X1 U174 ( .A1(n74), .A2(A_AND_B[12]), .ZN(A_XOR_B[12]) );
  NOR2_X1 U175 ( .A1(n75), .A2(A_AND_B[14]), .ZN(A_XOR_B[14]) );
  NOR2_X1 U176 ( .A1(n76), .A2(A_AND_B[15]), .ZN(A_XOR_B[15]) );
  NOR2_X1 U177 ( .A1(n77), .A2(A_AND_B[16]), .ZN(A_XOR_B[16]) );
  NOR2_X1 U178 ( .A1(n78), .A2(A_AND_B[17]), .ZN(A_XOR_B[17]) );
  NOR2_X1 U179 ( .A1(n79), .A2(A_AND_B[18]), .ZN(A_XOR_B[18]) );
  NOR2_X1 U180 ( .A1(n80), .A2(A_AND_B[19]), .ZN(A_XOR_B[19]) );
  NOR2_X1 U181 ( .A1(n81), .A2(A_AND_B[1]), .ZN(A_XOR_B[1]) );
  NOR2_X1 U182 ( .A1(n82), .A2(A_AND_B[20]), .ZN(A_XOR_B[20]) );
  NOR2_X1 U183 ( .A1(n83), .A2(A_AND_B[21]), .ZN(A_XOR_B[21]) );
  NOR2_X1 U184 ( .A1(n84), .A2(A_AND_B[22]), .ZN(A_XOR_B[22]) );
  NOR2_X1 U185 ( .A1(n85), .A2(A_AND_B[23]), .ZN(A_XOR_B[23]) );
  NOR2_X1 U186 ( .A1(n86), .A2(A_AND_B[24]), .ZN(A_XOR_B[24]) );
  NOR2_X1 U187 ( .A1(n87), .A2(A_AND_B[25]), .ZN(A_XOR_B[25]) );
  NOR2_X1 U188 ( .A1(n88), .A2(A_AND_B[26]), .ZN(A_XOR_B[26]) );
  NOR2_X1 U189 ( .A1(n89), .A2(A_AND_B[27]), .ZN(A_XOR_B[27]) );
  NOR2_X1 U190 ( .A1(n90), .A2(A_AND_B[28]), .ZN(A_XOR_B[28]) );
  NOR2_X1 U191 ( .A1(n91), .A2(A_AND_B[29]), .ZN(A_XOR_B[29]) );
  NOR2_X1 U192 ( .A1(n92), .A2(A_AND_B[2]), .ZN(A_XOR_B[2]) );
  NOR2_X1 U193 ( .A1(n94), .A2(A_AND_B[3]), .ZN(A_XOR_B[3]) );
  NOR2_X1 U194 ( .A1(n95), .A2(A_AND_B[4]), .ZN(A_XOR_B[4]) );
  NOR2_X1 U195 ( .A1(n96), .A2(A_AND_B[5]), .ZN(A_XOR_B[5]) );
  NOR2_X1 U196 ( .A1(n97), .A2(A_AND_B[6]), .ZN(A_XOR_B[6]) );
  NOR2_X1 U197 ( .A1(n98), .A2(A_AND_B[7]), .ZN(A_XOR_B[7]) );
  NOR2_X1 U198 ( .A1(n99), .A2(A_AND_B[8]), .ZN(A_XOR_B[8]) );
  NOR2_X1 U199 ( .A1(n100), .A2(A_AND_B[9]), .ZN(A_XOR_B[9]) );
endmodule


module ALU_N32 ( .FUNC({\FUNC[4] , \FUNC[3] , \FUNC[2] , \FUNC[1] , \FUNC[0] }
        ), DATA1, DATA2, OUT_ALU );
  input [31:0] DATA1;
  input [31:0] DATA2;
  output [31:0] OUT_ALU;
  input \FUNC[4] , \FUNC[3] , \FUNC[2] , \FUNC[1] , \FUNC[0] ;
  wire   add_sub, carry_out, \out_sgeu[0] , \out_sge[0] , \out_sgt[0] ,
         \out_sleu[0] , \out_sle[0] , \out_slt[0] , \out_sltu[0] ,
         \out_seq[0] , N121, N122, N123, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159;
  wire   [4:0] FUNC;
  wire   [31:0] out_barrel_shifter;
  wire   [31:0] out_st;
  wire   [31:0] out_not;
  wire   [31:0] out_and;
  wire   [31:0] out_xor;
  wire   [31:0] out_or;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106, SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        SYNOPSYS_UNCONNECTED__118, SYNOPSYS_UNCONNECTED__119, 
        SYNOPSYS_UNCONNECTED__120, SYNOPSYS_UNCONNECTED__121, 
        SYNOPSYS_UNCONNECTED__122, SYNOPSYS_UNCONNECTED__123, 
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        SYNOPSYS_UNCONNECTED__126, SYNOPSYS_UNCONNECTED__127, 
        SYNOPSYS_UNCONNECTED__128, SYNOPSYS_UNCONNECTED__129, 
        SYNOPSYS_UNCONNECTED__130, SYNOPSYS_UNCONNECTED__131, 
        SYNOPSYS_UNCONNECTED__132, SYNOPSYS_UNCONNECTED__133, 
        SYNOPSYS_UNCONNECTED__134, SYNOPSYS_UNCONNECTED__135, 
        SYNOPSYS_UNCONNECTED__136, SYNOPSYS_UNCONNECTED__137, 
        SYNOPSYS_UNCONNECTED__138, SYNOPSYS_UNCONNECTED__139, 
        SYNOPSYS_UNCONNECTED__140, SYNOPSYS_UNCONNECTED__141, 
        SYNOPSYS_UNCONNECTED__142, SYNOPSYS_UNCONNECTED__143, 
        SYNOPSYS_UNCONNECTED__144, SYNOPSYS_UNCONNECTED__145, 
        SYNOPSYS_UNCONNECTED__146, SYNOPSYS_UNCONNECTED__147, 
        SYNOPSYS_UNCONNECTED__148, SYNOPSYS_UNCONNECTED__149, 
        SYNOPSYS_UNCONNECTED__150, SYNOPSYS_UNCONNECTED__151, 
        SYNOPSYS_UNCONNECTED__152, SYNOPSYS_UNCONNECTED__153, 
        SYNOPSYS_UNCONNECTED__154, SYNOPSYS_UNCONNECTED__155, 
        SYNOPSYS_UNCONNECTED__156, SYNOPSYS_UNCONNECTED__157, 
        SYNOPSYS_UNCONNECTED__158, SYNOPSYS_UNCONNECTED__159, 
        SYNOPSYS_UNCONNECTED__160, SYNOPSYS_UNCONNECTED__161, 
        SYNOPSYS_UNCONNECTED__162, SYNOPSYS_UNCONNECTED__163, 
        SYNOPSYS_UNCONNECTED__164, SYNOPSYS_UNCONNECTED__165, 
        SYNOPSYS_UNCONNECTED__166, SYNOPSYS_UNCONNECTED__167, 
        SYNOPSYS_UNCONNECTED__168, SYNOPSYS_UNCONNECTED__169, 
        SYNOPSYS_UNCONNECTED__170, SYNOPSYS_UNCONNECTED__171, 
        SYNOPSYS_UNCONNECTED__172, SYNOPSYS_UNCONNECTED__173, 
        SYNOPSYS_UNCONNECTED__174, SYNOPSYS_UNCONNECTED__175, 
        SYNOPSYS_UNCONNECTED__176, SYNOPSYS_UNCONNECTED__177, 
        SYNOPSYS_UNCONNECTED__178, SYNOPSYS_UNCONNECTED__179, 
        SYNOPSYS_UNCONNECTED__180, SYNOPSYS_UNCONNECTED__181, 
        SYNOPSYS_UNCONNECTED__182, SYNOPSYS_UNCONNECTED__183, 
        SYNOPSYS_UNCONNECTED__184, SYNOPSYS_UNCONNECTED__185, 
        SYNOPSYS_UNCONNECTED__186, SYNOPSYS_UNCONNECTED__187, 
        SYNOPSYS_UNCONNECTED__188, SYNOPSYS_UNCONNECTED__189, 
        SYNOPSYS_UNCONNECTED__190, SYNOPSYS_UNCONNECTED__191, 
        SYNOPSYS_UNCONNECTED__192, SYNOPSYS_UNCONNECTED__193, 
        SYNOPSYS_UNCONNECTED__194, SYNOPSYS_UNCONNECTED__195, 
        SYNOPSYS_UNCONNECTED__196, SYNOPSYS_UNCONNECTED__197, 
        SYNOPSYS_UNCONNECTED__198, SYNOPSYS_UNCONNECTED__199, 
        SYNOPSYS_UNCONNECTED__200, SYNOPSYS_UNCONNECTED__201, 
        SYNOPSYS_UNCONNECTED__202, SYNOPSYS_UNCONNECTED__203, 
        SYNOPSYS_UNCONNECTED__204, SYNOPSYS_UNCONNECTED__205, 
        SYNOPSYS_UNCONNECTED__206, SYNOPSYS_UNCONNECTED__207, 
        SYNOPSYS_UNCONNECTED__208, SYNOPSYS_UNCONNECTED__209, 
        SYNOPSYS_UNCONNECTED__210, SYNOPSYS_UNCONNECTED__211, 
        SYNOPSYS_UNCONNECTED__212, SYNOPSYS_UNCONNECTED__213, 
        SYNOPSYS_UNCONNECTED__214, SYNOPSYS_UNCONNECTED__215, 
        SYNOPSYS_UNCONNECTED__216, SYNOPSYS_UNCONNECTED__217, 
        SYNOPSYS_UNCONNECTED__218, SYNOPSYS_UNCONNECTED__219, 
        SYNOPSYS_UNCONNECTED__220, SYNOPSYS_UNCONNECTED__221, 
        SYNOPSYS_UNCONNECTED__222, SYNOPSYS_UNCONNECTED__223, 
        SYNOPSYS_UNCONNECTED__224, SYNOPSYS_UNCONNECTED__225, 
        SYNOPSYS_UNCONNECTED__226, SYNOPSYS_UNCONNECTED__227, 
        SYNOPSYS_UNCONNECTED__228, SYNOPSYS_UNCONNECTED__229, 
        SYNOPSYS_UNCONNECTED__230, SYNOPSYS_UNCONNECTED__231, 
        SYNOPSYS_UNCONNECTED__232, SYNOPSYS_UNCONNECTED__233, 
        SYNOPSYS_UNCONNECTED__234, SYNOPSYS_UNCONNECTED__235, 
        SYNOPSYS_UNCONNECTED__236, SYNOPSYS_UNCONNECTED__237, 
        SYNOPSYS_UNCONNECTED__238, SYNOPSYS_UNCONNECTED__239, 
        SYNOPSYS_UNCONNECTED__240, SYNOPSYS_UNCONNECTED__241, 
        SYNOPSYS_UNCONNECTED__242, SYNOPSYS_UNCONNECTED__243, 
        SYNOPSYS_UNCONNECTED__244, SYNOPSYS_UNCONNECTED__245, 
        SYNOPSYS_UNCONNECTED__246, SYNOPSYS_UNCONNECTED__247;

  barrel_shifter_Nbit32 BRRL_SHFT ( .A(DATA1), .B({DATA2[31:3], n24, DATA2[1], 
        n20}), .SHIFT_ROTATE(N121), .LOGIC_ARITH(N122), .LEFT_RIGHT(N123), 
        .OUTPUT(out_barrel_shifter) );
  ADDER_P4_N_BIT32_1 SPARSE_TREE_ADDER ( .A(DATA1), .B(DATA2), .add_sub(
        add_sub), .Cout(carry_out), .SUM(out_st) );
  LOGIC_BLOCK_N32 LGC_BLOCK ( .SUM(out_st), .C_OUT(carry_out), .A(DATA1), .B({
        DATA2[31:3], n24, DATA2[1], n20}), .A_GEU_B({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, SYNOPSYS_UNCONNECTED__22, 
        SYNOPSYS_UNCONNECTED__23, SYNOPSYS_UNCONNECTED__24, 
        SYNOPSYS_UNCONNECTED__25, SYNOPSYS_UNCONNECTED__26, 
        SYNOPSYS_UNCONNECTED__27, SYNOPSYS_UNCONNECTED__28, 
        SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, \out_sgeu[0] }), 
        .A_GE_B({SYNOPSYS_UNCONNECTED__31, SYNOPSYS_UNCONNECTED__32, 
        SYNOPSYS_UNCONNECTED__33, SYNOPSYS_UNCONNECTED__34, 
        SYNOPSYS_UNCONNECTED__35, SYNOPSYS_UNCONNECTED__36, 
        SYNOPSYS_UNCONNECTED__37, SYNOPSYS_UNCONNECTED__38, 
        SYNOPSYS_UNCONNECTED__39, SYNOPSYS_UNCONNECTED__40, 
        SYNOPSYS_UNCONNECTED__41, SYNOPSYS_UNCONNECTED__42, 
        SYNOPSYS_UNCONNECTED__43, SYNOPSYS_UNCONNECTED__44, 
        SYNOPSYS_UNCONNECTED__45, SYNOPSYS_UNCONNECTED__46, 
        SYNOPSYS_UNCONNECTED__47, SYNOPSYS_UNCONNECTED__48, 
        SYNOPSYS_UNCONNECTED__49, SYNOPSYS_UNCONNECTED__50, 
        SYNOPSYS_UNCONNECTED__51, SYNOPSYS_UNCONNECTED__52, 
        SYNOPSYS_UNCONNECTED__53, SYNOPSYS_UNCONNECTED__54, 
        SYNOPSYS_UNCONNECTED__55, SYNOPSYS_UNCONNECTED__56, 
        SYNOPSYS_UNCONNECTED__57, SYNOPSYS_UNCONNECTED__58, 
        SYNOPSYS_UNCONNECTED__59, SYNOPSYS_UNCONNECTED__60, 
        SYNOPSYS_UNCONNECTED__61, \out_sge[0] }), .A_GT_B({
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, \out_sgt[0] }), .A_LEU_B({
        SYNOPSYS_UNCONNECTED__93, SYNOPSYS_UNCONNECTED__94, 
        SYNOPSYS_UNCONNECTED__95, SYNOPSYS_UNCONNECTED__96, 
        SYNOPSYS_UNCONNECTED__97, SYNOPSYS_UNCONNECTED__98, 
        SYNOPSYS_UNCONNECTED__99, SYNOPSYS_UNCONNECTED__100, 
        SYNOPSYS_UNCONNECTED__101, SYNOPSYS_UNCONNECTED__102, 
        SYNOPSYS_UNCONNECTED__103, SYNOPSYS_UNCONNECTED__104, 
        SYNOPSYS_UNCONNECTED__105, SYNOPSYS_UNCONNECTED__106, 
        SYNOPSYS_UNCONNECTED__107, SYNOPSYS_UNCONNECTED__108, 
        SYNOPSYS_UNCONNECTED__109, SYNOPSYS_UNCONNECTED__110, 
        SYNOPSYS_UNCONNECTED__111, SYNOPSYS_UNCONNECTED__112, 
        SYNOPSYS_UNCONNECTED__113, SYNOPSYS_UNCONNECTED__114, 
        SYNOPSYS_UNCONNECTED__115, SYNOPSYS_UNCONNECTED__116, 
        SYNOPSYS_UNCONNECTED__117, SYNOPSYS_UNCONNECTED__118, 
        SYNOPSYS_UNCONNECTED__119, SYNOPSYS_UNCONNECTED__120, 
        SYNOPSYS_UNCONNECTED__121, SYNOPSYS_UNCONNECTED__122, 
        SYNOPSYS_UNCONNECTED__123, \out_sleu[0] }), .A_LE_B({
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        SYNOPSYS_UNCONNECTED__126, SYNOPSYS_UNCONNECTED__127, 
        SYNOPSYS_UNCONNECTED__128, SYNOPSYS_UNCONNECTED__129, 
        SYNOPSYS_UNCONNECTED__130, SYNOPSYS_UNCONNECTED__131, 
        SYNOPSYS_UNCONNECTED__132, SYNOPSYS_UNCONNECTED__133, 
        SYNOPSYS_UNCONNECTED__134, SYNOPSYS_UNCONNECTED__135, 
        SYNOPSYS_UNCONNECTED__136, SYNOPSYS_UNCONNECTED__137, 
        SYNOPSYS_UNCONNECTED__138, SYNOPSYS_UNCONNECTED__139, 
        SYNOPSYS_UNCONNECTED__140, SYNOPSYS_UNCONNECTED__141, 
        SYNOPSYS_UNCONNECTED__142, SYNOPSYS_UNCONNECTED__143, 
        SYNOPSYS_UNCONNECTED__144, SYNOPSYS_UNCONNECTED__145, 
        SYNOPSYS_UNCONNECTED__146, SYNOPSYS_UNCONNECTED__147, 
        SYNOPSYS_UNCONNECTED__148, SYNOPSYS_UNCONNECTED__149, 
        SYNOPSYS_UNCONNECTED__150, SYNOPSYS_UNCONNECTED__151, 
        SYNOPSYS_UNCONNECTED__152, SYNOPSYS_UNCONNECTED__153, 
        SYNOPSYS_UNCONNECTED__154, \out_sle[0] }), .A_LT_B({
        SYNOPSYS_UNCONNECTED__155, SYNOPSYS_UNCONNECTED__156, 
        SYNOPSYS_UNCONNECTED__157, SYNOPSYS_UNCONNECTED__158, 
        SYNOPSYS_UNCONNECTED__159, SYNOPSYS_UNCONNECTED__160, 
        SYNOPSYS_UNCONNECTED__161, SYNOPSYS_UNCONNECTED__162, 
        SYNOPSYS_UNCONNECTED__163, SYNOPSYS_UNCONNECTED__164, 
        SYNOPSYS_UNCONNECTED__165, SYNOPSYS_UNCONNECTED__166, 
        SYNOPSYS_UNCONNECTED__167, SYNOPSYS_UNCONNECTED__168, 
        SYNOPSYS_UNCONNECTED__169, SYNOPSYS_UNCONNECTED__170, 
        SYNOPSYS_UNCONNECTED__171, SYNOPSYS_UNCONNECTED__172, 
        SYNOPSYS_UNCONNECTED__173, SYNOPSYS_UNCONNECTED__174, 
        SYNOPSYS_UNCONNECTED__175, SYNOPSYS_UNCONNECTED__176, 
        SYNOPSYS_UNCONNECTED__177, SYNOPSYS_UNCONNECTED__178, 
        SYNOPSYS_UNCONNECTED__179, SYNOPSYS_UNCONNECTED__180, 
        SYNOPSYS_UNCONNECTED__181, SYNOPSYS_UNCONNECTED__182, 
        SYNOPSYS_UNCONNECTED__183, SYNOPSYS_UNCONNECTED__184, 
        SYNOPSYS_UNCONNECTED__185, \out_slt[0] }), .A_LTU_B({
        SYNOPSYS_UNCONNECTED__186, SYNOPSYS_UNCONNECTED__187, 
        SYNOPSYS_UNCONNECTED__188, SYNOPSYS_UNCONNECTED__189, 
        SYNOPSYS_UNCONNECTED__190, SYNOPSYS_UNCONNECTED__191, 
        SYNOPSYS_UNCONNECTED__192, SYNOPSYS_UNCONNECTED__193, 
        SYNOPSYS_UNCONNECTED__194, SYNOPSYS_UNCONNECTED__195, 
        SYNOPSYS_UNCONNECTED__196, SYNOPSYS_UNCONNECTED__197, 
        SYNOPSYS_UNCONNECTED__198, SYNOPSYS_UNCONNECTED__199, 
        SYNOPSYS_UNCONNECTED__200, SYNOPSYS_UNCONNECTED__201, 
        SYNOPSYS_UNCONNECTED__202, SYNOPSYS_UNCONNECTED__203, 
        SYNOPSYS_UNCONNECTED__204, SYNOPSYS_UNCONNECTED__205, 
        SYNOPSYS_UNCONNECTED__206, SYNOPSYS_UNCONNECTED__207, 
        SYNOPSYS_UNCONNECTED__208, SYNOPSYS_UNCONNECTED__209, 
        SYNOPSYS_UNCONNECTED__210, SYNOPSYS_UNCONNECTED__211, 
        SYNOPSYS_UNCONNECTED__212, SYNOPSYS_UNCONNECTED__213, 
        SYNOPSYS_UNCONNECTED__214, SYNOPSYS_UNCONNECTED__215, 
        SYNOPSYS_UNCONNECTED__216, \out_sltu[0] }), .A_EQ_B({
        SYNOPSYS_UNCONNECTED__217, SYNOPSYS_UNCONNECTED__218, 
        SYNOPSYS_UNCONNECTED__219, SYNOPSYS_UNCONNECTED__220, 
        SYNOPSYS_UNCONNECTED__221, SYNOPSYS_UNCONNECTED__222, 
        SYNOPSYS_UNCONNECTED__223, SYNOPSYS_UNCONNECTED__224, 
        SYNOPSYS_UNCONNECTED__225, SYNOPSYS_UNCONNECTED__226, 
        SYNOPSYS_UNCONNECTED__227, SYNOPSYS_UNCONNECTED__228, 
        SYNOPSYS_UNCONNECTED__229, SYNOPSYS_UNCONNECTED__230, 
        SYNOPSYS_UNCONNECTED__231, SYNOPSYS_UNCONNECTED__232, 
        SYNOPSYS_UNCONNECTED__233, SYNOPSYS_UNCONNECTED__234, 
        SYNOPSYS_UNCONNECTED__235, SYNOPSYS_UNCONNECTED__236, 
        SYNOPSYS_UNCONNECTED__237, SYNOPSYS_UNCONNECTED__238, 
        SYNOPSYS_UNCONNECTED__239, SYNOPSYS_UNCONNECTED__240, 
        SYNOPSYS_UNCONNECTED__241, SYNOPSYS_UNCONNECTED__242, 
        SYNOPSYS_UNCONNECTED__243, SYNOPSYS_UNCONNECTED__244, 
        SYNOPSYS_UNCONNECTED__245, SYNOPSYS_UNCONNECTED__246, 
        SYNOPSYS_UNCONNECTED__247, \out_seq[0] }), .NOT_A(out_not), .A_AND_B(
        out_and), .A_XOR_B(out_xor), .A_OR_B(out_or) );
  INV_X1 U3 ( .A(n51), .ZN(n9) );
  AOI22_X1 U4 ( .A1(out_or[9]), .A2(n28), .B1(n56), .B2(out_xor[9]), .ZN(n1)
         );
  NAND3_X1 U5 ( .A1(n158), .A2(n159), .A3(n1), .ZN(OUT_ALU[9]) );
  AOI22_X1 U6 ( .A1(out_st[13]), .A2(n65), .B1(n157), .B2(
        out_barrel_shifter[13]), .ZN(n2) );
  AOI22_X1 U7 ( .A1(out_not[13]), .A2(n45), .B1(out_and[13]), .B2(n67), .ZN(n3) );
  AOI22_X1 U8 ( .A1(out_or[13]), .A2(n43), .B1(n42), .B2(out_xor[13]), .ZN(n4)
         );
  NAND3_X1 U9 ( .A1(n2), .A2(n3), .A3(n4), .ZN(OUT_ALU[13]) );
  AOI22_X1 U10 ( .A1(out_st[30]), .A2(n44), .B1(n46), .B2(
        out_barrel_shifter[30]), .ZN(n5) );
  AOI22_X1 U11 ( .A1(out_not[30]), .A2(n45), .B1(out_and[30]), .B2(n67), .ZN(
        n6) );
  AOI22_X1 U12 ( .A1(out_or[30]), .A2(n28), .B1(n56), .B2(out_xor[30]), .ZN(n7) );
  NAND3_X1 U13 ( .A1(n5), .A2(n6), .A3(n7), .ZN(OUT_ALU[30]) );
  AOI22_X1 U14 ( .A1(out_not[18]), .A2(n66), .B1(out_and[18]), .B2(n67), .ZN(
        n8) );
  NAND3_X1 U15 ( .A1(n95), .A2(n96), .A3(n8), .ZN(OUT_ALU[18]) );
  AND2_X1 U16 ( .A1(\out_sgt[0] ), .A2(n9), .ZN(n31) );
  CLKBUF_X1 U17 ( .A(DATA2[0]), .Z(n20) );
  INV_X1 U18 ( .A(n71), .ZN(n10) );
  NOR2_X2 U19 ( .A1(n73), .A2(n68), .ZN(N122) );
  BUF_X1 U20 ( .A(n10), .Z(n25) );
  NOR3_X2 U21 ( .A1(n51), .A2(n11), .A3(n52), .ZN(n66) );
  INV_X1 U22 ( .A(n68), .ZN(n11) );
  OAI21_X1 U23 ( .B1(n68), .B2(n71), .A(FUNC[1]), .ZN(N123) );
  BUF_X1 U24 ( .A(DATA2[2]), .Z(n24) );
  INV_X1 U25 ( .A(FUNC[2]), .ZN(n52) );
  AND2_X2 U26 ( .A1(n50), .A2(n73), .ZN(n67) );
  BUF_X1 U27 ( .A(n65), .Z(n44) );
  BUF_X1 U28 ( .A(n157), .Z(n46) );
  BUF_X1 U29 ( .A(n56), .Z(n42) );
  BUF_X1 U30 ( .A(n66), .Z(n45) );
  AND2_X1 U31 ( .A1(n40), .A2(FUNC[0]), .ZN(n27) );
  NAND2_X1 U32 ( .A1(n81), .A2(n21), .ZN(OUT_ALU[12]) );
  NOR2_X1 U33 ( .A1(n23), .A2(n22), .ZN(n21) );
  INV_X1 U34 ( .A(n82), .ZN(n22) );
  INV_X1 U35 ( .A(n80), .ZN(n23) );
  NAND2_X1 U36 ( .A1(\out_sle[0] ), .A2(n26), .ZN(n55) );
  AND2_X1 U37 ( .A1(n52), .A2(n73), .ZN(n26) );
  NAND3_X1 U38 ( .A1(n27), .A2(n41), .A3(n39), .ZN(add_sub) );
  NOR2_X2 U39 ( .A1(n49), .A2(n53), .ZN(n56) );
  INV_X1 U40 ( .A(FUNC[1]), .ZN(n69) );
  INV_X1 U41 ( .A(FUNC[3]), .ZN(n68) );
  NOR2_X2 U42 ( .A1(n49), .A2(n47), .ZN(n65) );
  INV_X1 U43 ( .A(FUNC[1]), .ZN(n39) );
  INV_X1 U44 ( .A(FUNC[4]), .ZN(n40) );
  NOR2_X1 U45 ( .A1(FUNC[3]), .A2(FUNC[2]), .ZN(n41) );
  INV_X1 U46 ( .A(FUNC[0]), .ZN(n71) );
  OAI21_X2 U47 ( .B1(n53), .B2(n70), .A(n48), .ZN(n157) );
  AOI22_X1 U48 ( .A1(out_xor[14]), .A2(n42), .B1(n43), .B2(out_or[14]), .ZN(
        n83) );
  AOI22_X1 U49 ( .A1(out_xor[3]), .A2(n42), .B1(n28), .B2(out_or[3]), .ZN(n139) );
  AOI22_X1 U50 ( .A1(out_xor[12]), .A2(n42), .B1(n43), .B2(out_or[12]), .ZN(
        n80) );
  AOI22_X1 U51 ( .A1(out_xor[11]), .A2(n42), .B1(n28), .B2(out_or[11]), .ZN(
        n77) );
  AOI22_X1 U52 ( .A1(out_xor[7]), .A2(n56), .B1(n28), .B2(out_or[7]), .ZN(n151) );
  AOI22_X1 U53 ( .A1(out_xor[10]), .A2(n42), .B1(n28), .B2(out_or[10]), .ZN(
        n74) );
  AOI22_X1 U54 ( .A1(out_xor[18]), .A2(n42), .B1(n28), .B2(out_or[18]), .ZN(
        n95) );
  AOI22_X1 U55 ( .A1(out_xor[17]), .A2(n42), .B1(n43), .B2(out_or[17]), .ZN(
        n92) );
  AOI22_X1 U56 ( .A1(out_xor[15]), .A2(n42), .B1(n43), .B2(out_or[15]), .ZN(
        n86) );
  AOI22_X1 U57 ( .A1(out_xor[25]), .A2(n56), .B1(n28), .B2(out_or[25]), .ZN(
        n118) );
  AOI22_X1 U58 ( .A1(out_xor[24]), .A2(n42), .B1(n28), .B2(out_or[24]), .ZN(
        n115) );
  AOI22_X1 U59 ( .A1(out_xor[23]), .A2(n56), .B1(n28), .B2(out_or[23]), .ZN(
        n112) );
  AOI22_X1 U60 ( .A1(out_xor[22]), .A2(n56), .B1(n28), .B2(out_or[22]), .ZN(
        n109) );
  AOI22_X1 U61 ( .A1(out_xor[29]), .A2(n56), .B1(n28), .B2(out_or[29]), .ZN(
        n130) );
  AOI22_X1 U62 ( .A1(out_xor[28]), .A2(n42), .B1(n28), .B2(out_or[28]), .ZN(
        n127) );
  AOI22_X1 U63 ( .A1(out_xor[27]), .A2(n56), .B1(n28), .B2(out_or[27]), .ZN(
        n124) );
  AOI22_X1 U64 ( .A1(out_xor[26]), .A2(n56), .B1(n28), .B2(out_or[26]), .ZN(
        n121) );
  AOI22_X1 U65 ( .A1(out_xor[21]), .A2(n56), .B1(n28), .B2(out_or[21]), .ZN(
        n106) );
  AOI22_X1 U66 ( .A1(out_xor[20]), .A2(n42), .B1(n28), .B2(out_or[20]), .ZN(
        n103) );
  AOI22_X1 U67 ( .A1(out_xor[1]), .A2(n42), .B1(n28), .B2(out_or[1]), .ZN(n100) );
  AOI22_X1 U68 ( .A1(out_xor[19]), .A2(n42), .B1(n28), .B2(out_or[19]), .ZN(
        n97) );
  AOI22_X1 U69 ( .A1(out_xor[2]), .A2(n56), .B1(n28), .B2(out_or[2]), .ZN(n133) );
  AOI22_X1 U70 ( .A1(out_xor[31]), .A2(n56), .B1(out_or[31]), .B2(n43), .ZN(
        n136) );
  AOI22_X1 U71 ( .A1(out_xor[8]), .A2(n42), .B1(n28), .B2(out_or[8]), .ZN(n154) );
  AOI22_X1 U72 ( .A1(out_xor[6]), .A2(n42), .B1(n28), .B2(out_or[6]), .ZN(n148) );
  AOI22_X1 U73 ( .A1(out_xor[5]), .A2(n42), .B1(n28), .B2(out_or[5]), .ZN(n145) );
  AOI22_X1 U74 ( .A1(out_xor[4]), .A2(n42), .B1(n28), .B2(out_or[4]), .ZN(n142) );
  AOI21_X1 U75 ( .B1(out_barrel_shifter[0]), .B2(n157), .A(n61), .ZN(n62) );
  NAND4_X1 U76 ( .A1(n60), .A2(n59), .A3(n58), .A4(n57), .ZN(n61) );
  NAND2_X1 U77 ( .A1(out_or[0]), .A2(n43), .ZN(n57) );
  NAND2_X1 U78 ( .A1(out_xor[0]), .A2(n42), .ZN(n58) );
  AOI22_X1 U79 ( .A1(out_and[0]), .A2(n67), .B1(n45), .B2(out_not[0]), .ZN(n59) );
  NAND2_X1 U80 ( .A1(out_st[0]), .A2(n44), .ZN(n60) );
  NAND2_X1 U81 ( .A1(n71), .A2(n30), .ZN(n29) );
  INV_X1 U82 ( .A(n52), .ZN(n30) );
  OAI21_X1 U83 ( .B1(\out_seq[0] ), .B2(n52), .A(n25), .ZN(n35) );
  AOI22_X1 U84 ( .A1(out_xor[16]), .A2(n42), .B1(n43), .B2(out_or[16]), .ZN(
        n89) );
  BUF_X1 U85 ( .A(n28), .Z(n43) );
  NAND2_X1 U86 ( .A1(n52), .A2(n11), .ZN(n48) );
  INV_X1 U87 ( .A(n53), .ZN(n47) );
  NAND2_X1 U88 ( .A1(n50), .A2(n52), .ZN(n49) );
  NAND2_X1 U89 ( .A1(n71), .A2(FUNC[1]), .ZN(n51) );
  NOR2_X1 U90 ( .A1(FUNC[4]), .A2(FUNC[3]), .ZN(n50) );
  AND4_X1 U91 ( .A1(n50), .A2(n25), .A3(FUNC[2]), .A4(n69), .ZN(n28) );
  OR2_X1 U92 ( .A1(\out_seq[0] ), .A2(n29), .ZN(n38) );
  OAI21_X1 U93 ( .B1(n32), .B2(n31), .A(n30), .ZN(n54) );
  OAI21_X1 U94 ( .B1(\out_sleu[0] ), .B2(n53), .A(n72), .ZN(n32) );
  OAI211_X1 U95 ( .C1(n35), .C2(n36), .A(n38), .B(n33), .ZN(n37) );
  NAND2_X1 U96 ( .A1(\out_sltu[0] ), .A2(n34), .ZN(n33) );
  NOR2_X1 U97 ( .A1(n71), .A2(n69), .ZN(n34) );
  AOI21_X1 U98 ( .B1(\out_sleu[0] ), .B2(n69), .A(FUNC[2]), .ZN(n36) );
  AOI21_X1 U99 ( .B1(\out_slt[0] ), .B2(n9), .A(n37), .ZN(n64) );
  NAND2_X1 U100 ( .A1(n25), .A2(FUNC[1]), .ZN(n53) );
  OAI211_X1 U101 ( .C1(n64), .C2(n40), .A(n63), .B(n62), .ZN(OUT_ALU[0]) );
  MUX2_X1 U102 ( .A(n55), .B(n54), .S(n11), .Z(n63) );
  NOR2_X1 U103 ( .A1(FUNC[2]), .A2(n69), .ZN(N121) );
  NOR2_X1 U104 ( .A1(n10), .A2(FUNC[1]), .ZN(n73) );
  NAND2_X1 U105 ( .A1(n30), .A2(n68), .ZN(n70) );
  OAI221_X1 U106 ( .B1(n25), .B2(\out_sge[0] ), .C1(n71), .C2(\out_sgeu[0] ), 
        .A(n69), .ZN(n72) );
  AOI22_X1 U107 ( .A1(n67), .A2(out_and[10]), .B1(n45), .B2(out_not[10]), .ZN(
        n76) );
  AOI22_X1 U108 ( .A1(out_st[10]), .A2(n44), .B1(out_barrel_shifter[10]), .B2(
        n46), .ZN(n75) );
  NAND3_X1 U109 ( .A1(n75), .A2(n76), .A3(n74), .ZN(OUT_ALU[10]) );
  AOI22_X1 U110 ( .A1(n67), .A2(out_and[11]), .B1(n66), .B2(out_not[11]), .ZN(
        n79) );
  AOI22_X1 U111 ( .A1(out_st[11]), .A2(n65), .B1(out_barrel_shifter[11]), .B2(
        n157), .ZN(n78) );
  NAND3_X1 U112 ( .A1(n79), .A2(n78), .A3(n77), .ZN(OUT_ALU[11]) );
  AOI22_X1 U113 ( .A1(n67), .A2(out_and[12]), .B1(n66), .B2(out_not[12]), .ZN(
        n82) );
  AOI22_X1 U114 ( .A1(out_st[12]), .A2(n65), .B1(out_barrel_shifter[12]), .B2(
        n157), .ZN(n81) );
  AOI22_X1 U115 ( .A1(n67), .A2(out_and[14]), .B1(n66), .B2(out_not[14]), .ZN(
        n85) );
  AOI22_X1 U116 ( .A1(out_st[14]), .A2(n65), .B1(out_barrel_shifter[14]), .B2(
        n157), .ZN(n84) );
  NAND3_X1 U117 ( .A1(n85), .A2(n84), .A3(n83), .ZN(OUT_ALU[14]) );
  AOI22_X1 U118 ( .A1(n67), .A2(out_and[15]), .B1(n66), .B2(out_not[15]), .ZN(
        n88) );
  AOI22_X1 U119 ( .A1(out_st[15]), .A2(n65), .B1(out_barrel_shifter[15]), .B2(
        n157), .ZN(n87) );
  NAND3_X1 U120 ( .A1(n88), .A2(n87), .A3(n86), .ZN(OUT_ALU[15]) );
  AOI22_X1 U121 ( .A1(n67), .A2(out_and[16]), .B1(n66), .B2(out_not[16]), .ZN(
        n91) );
  AOI22_X1 U122 ( .A1(out_st[16]), .A2(n65), .B1(out_barrel_shifter[16]), .B2(
        n157), .ZN(n90) );
  NAND3_X1 U123 ( .A1(n90), .A2(n91), .A3(n89), .ZN(OUT_ALU[16]) );
  AOI22_X1 U124 ( .A1(n67), .A2(out_and[17]), .B1(n66), .B2(out_not[17]), .ZN(
        n94) );
  AOI22_X1 U125 ( .A1(out_st[17]), .A2(n65), .B1(out_barrel_shifter[17]), .B2(
        n157), .ZN(n93) );
  NAND3_X1 U126 ( .A1(n94), .A2(n93), .A3(n92), .ZN(OUT_ALU[17]) );
  AOI22_X1 U127 ( .A1(out_st[18]), .A2(n65), .B1(out_barrel_shifter[18]), .B2(
        n157), .ZN(n96) );
  AOI22_X1 U128 ( .A1(n67), .A2(out_and[19]), .B1(n45), .B2(out_not[19]), .ZN(
        n99) );
  AOI22_X1 U129 ( .A1(out_st[19]), .A2(n65), .B1(out_barrel_shifter[19]), .B2(
        n157), .ZN(n98) );
  NAND3_X1 U130 ( .A1(n99), .A2(n98), .A3(n97), .ZN(OUT_ALU[19]) );
  AOI22_X1 U131 ( .A1(n67), .A2(out_and[1]), .B1(n66), .B2(out_not[1]), .ZN(
        n102) );
  AOI22_X1 U132 ( .A1(out_st[1]), .A2(n65), .B1(out_barrel_shifter[1]), .B2(
        n157), .ZN(n101) );
  NAND3_X1 U133 ( .A1(n102), .A2(n101), .A3(n100), .ZN(OUT_ALU[1]) );
  AOI22_X1 U134 ( .A1(n67), .A2(out_and[20]), .B1(n66), .B2(out_not[20]), .ZN(
        n105) );
  AOI22_X1 U135 ( .A1(out_st[20]), .A2(n65), .B1(out_barrel_shifter[20]), .B2(
        n157), .ZN(n104) );
  NAND3_X1 U136 ( .A1(n105), .A2(n104), .A3(n103), .ZN(OUT_ALU[20]) );
  AOI22_X1 U137 ( .A1(n67), .A2(out_and[21]), .B1(n66), .B2(out_not[21]), .ZN(
        n108) );
  AOI22_X1 U138 ( .A1(out_st[21]), .A2(n65), .B1(out_barrel_shifter[21]), .B2(
        n157), .ZN(n107) );
  NAND3_X1 U139 ( .A1(n108), .A2(n107), .A3(n106), .ZN(OUT_ALU[21]) );
  AOI22_X1 U140 ( .A1(n67), .A2(out_and[22]), .B1(n66), .B2(out_not[22]), .ZN(
        n111) );
  AOI22_X1 U141 ( .A1(out_st[22]), .A2(n65), .B1(out_barrel_shifter[22]), .B2(
        n157), .ZN(n110) );
  NAND3_X1 U142 ( .A1(n111), .A2(n110), .A3(n109), .ZN(OUT_ALU[22]) );
  AOI22_X1 U143 ( .A1(n67), .A2(out_and[23]), .B1(n66), .B2(out_not[23]), .ZN(
        n114) );
  AOI22_X1 U144 ( .A1(out_st[23]), .A2(n44), .B1(out_barrel_shifter[23]), .B2(
        n157), .ZN(n113) );
  NAND3_X1 U145 ( .A1(n114), .A2(n113), .A3(n112), .ZN(OUT_ALU[23]) );
  AOI22_X1 U146 ( .A1(n67), .A2(out_and[24]), .B1(n45), .B2(out_not[24]), .ZN(
        n117) );
  AOI22_X1 U147 ( .A1(out_st[24]), .A2(n44), .B1(out_barrel_shifter[24]), .B2(
        n157), .ZN(n116) );
  NAND3_X1 U148 ( .A1(n117), .A2(n116), .A3(n115), .ZN(OUT_ALU[24]) );
  AOI22_X1 U149 ( .A1(n67), .A2(out_and[25]), .B1(n45), .B2(out_not[25]), .ZN(
        n120) );
  AOI22_X1 U150 ( .A1(out_st[25]), .A2(n44), .B1(out_barrel_shifter[25]), .B2(
        n157), .ZN(n119) );
  NAND3_X1 U151 ( .A1(n120), .A2(n119), .A3(n118), .ZN(OUT_ALU[25]) );
  AOI22_X1 U152 ( .A1(n67), .A2(out_and[26]), .B1(n45), .B2(out_not[26]), .ZN(
        n123) );
  AOI22_X1 U153 ( .A1(out_st[26]), .A2(n44), .B1(out_barrel_shifter[26]), .B2(
        n157), .ZN(n122) );
  NAND3_X1 U154 ( .A1(n123), .A2(n122), .A3(n121), .ZN(OUT_ALU[26]) );
  AOI22_X1 U155 ( .A1(n67), .A2(out_and[27]), .B1(n45), .B2(out_not[27]), .ZN(
        n126) );
  AOI22_X1 U156 ( .A1(out_st[27]), .A2(n44), .B1(out_barrel_shifter[27]), .B2(
        n46), .ZN(n125) );
  NAND3_X1 U157 ( .A1(n126), .A2(n125), .A3(n124), .ZN(OUT_ALU[27]) );
  AOI22_X1 U158 ( .A1(n67), .A2(out_and[28]), .B1(n45), .B2(out_not[28]), .ZN(
        n129) );
  AOI22_X1 U159 ( .A1(out_st[28]), .A2(n44), .B1(out_barrel_shifter[28]), .B2(
        n46), .ZN(n128) );
  NAND3_X1 U160 ( .A1(n129), .A2(n128), .A3(n127), .ZN(OUT_ALU[28]) );
  AOI22_X1 U161 ( .A1(n67), .A2(out_and[29]), .B1(n45), .B2(out_not[29]), .ZN(
        n132) );
  AOI22_X1 U162 ( .A1(out_st[29]), .A2(n44), .B1(out_barrel_shifter[29]), .B2(
        n46), .ZN(n131) );
  NAND3_X1 U163 ( .A1(n132), .A2(n131), .A3(n130), .ZN(OUT_ALU[29]) );
  AOI22_X1 U164 ( .A1(n67), .A2(out_and[2]), .B1(n45), .B2(out_not[2]), .ZN(
        n135) );
  AOI22_X1 U165 ( .A1(out_st[2]), .A2(n44), .B1(out_barrel_shifter[2]), .B2(
        n46), .ZN(n134) );
  NAND3_X1 U166 ( .A1(n135), .A2(n134), .A3(n133), .ZN(OUT_ALU[2]) );
  AOI22_X1 U167 ( .A1(n67), .A2(out_and[31]), .B1(n45), .B2(out_not[31]), .ZN(
        n138) );
  AOI22_X1 U168 ( .A1(out_st[31]), .A2(n44), .B1(out_barrel_shifter[31]), .B2(
        n46), .ZN(n137) );
  NAND3_X1 U169 ( .A1(n138), .A2(n137), .A3(n136), .ZN(OUT_ALU[31]) );
  AOI22_X1 U170 ( .A1(n67), .A2(out_and[3]), .B1(n45), .B2(out_not[3]), .ZN(
        n141) );
  AOI22_X1 U171 ( .A1(out_st[3]), .A2(n44), .B1(out_barrel_shifter[3]), .B2(
        n46), .ZN(n140) );
  NAND3_X1 U172 ( .A1(n141), .A2(n140), .A3(n139), .ZN(OUT_ALU[3]) );
  AOI22_X1 U173 ( .A1(n67), .A2(out_and[4]), .B1(n45), .B2(out_not[4]), .ZN(
        n144) );
  AOI22_X1 U174 ( .A1(out_st[4]), .A2(n44), .B1(out_barrel_shifter[4]), .B2(
        n46), .ZN(n143) );
  NAND3_X1 U175 ( .A1(n144), .A2(n143), .A3(n142), .ZN(OUT_ALU[4]) );
  AOI22_X1 U176 ( .A1(n67), .A2(out_and[5]), .B1(n45), .B2(out_not[5]), .ZN(
        n147) );
  AOI22_X1 U177 ( .A1(out_st[5]), .A2(n44), .B1(out_barrel_shifter[5]), .B2(
        n46), .ZN(n146) );
  NAND3_X1 U178 ( .A1(n147), .A2(n146), .A3(n145), .ZN(OUT_ALU[5]) );
  AOI22_X1 U179 ( .A1(n67), .A2(out_and[6]), .B1(n45), .B2(out_not[6]), .ZN(
        n150) );
  AOI22_X1 U180 ( .A1(out_st[6]), .A2(n44), .B1(out_barrel_shifter[6]), .B2(
        n46), .ZN(n149) );
  NAND3_X1 U181 ( .A1(n150), .A2(n149), .A3(n148), .ZN(OUT_ALU[6]) );
  AOI22_X1 U182 ( .A1(n67), .A2(out_and[7]), .B1(n45), .B2(out_not[7]), .ZN(
        n153) );
  AOI22_X1 U183 ( .A1(out_st[7]), .A2(n44), .B1(out_barrel_shifter[7]), .B2(
        n46), .ZN(n152) );
  NAND3_X1 U184 ( .A1(n153), .A2(n152), .A3(n151), .ZN(OUT_ALU[7]) );
  AOI22_X1 U185 ( .A1(n67), .A2(out_and[8]), .B1(n45), .B2(out_not[8]), .ZN(
        n156) );
  AOI22_X1 U186 ( .A1(out_st[8]), .A2(n44), .B1(out_barrel_shifter[8]), .B2(
        n46), .ZN(n155) );
  NAND3_X1 U187 ( .A1(n156), .A2(n155), .A3(n154), .ZN(OUT_ALU[8]) );
  AOI22_X1 U188 ( .A1(n67), .A2(out_and[9]), .B1(n45), .B2(out_not[9]), .ZN(
        n159) );
  AOI22_X1 U189 ( .A1(out_st[9]), .A2(n44), .B1(out_barrel_shifter[9]), .B2(
        n46), .ZN(n158) );
endmodule


module PG_NETWORK_958 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_957 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op1), .A2(op2), .ZN(g) );
  XOR2_X1 U2 ( .A(op1), .B(op2), .Z(p) );
endmodule


module PG_NETWORK_956 ( op1, op2, g, p );
  input op1, op2;
  output g, p;
  wire   n1;

  XNOR2_X1 U1 ( .A(op1), .B(n1), .ZN(p) );
  INV_X1 U2 ( .A(op2), .ZN(n1) );
  AND2_X1 U3 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_955 ( op1, op2, g, p );
  input op1, op2;
  output g, p;
  wire   n1;

  XNOR2_X1 U1 ( .A(op1), .B(n1), .ZN(p) );
  INV_X1 U2 ( .A(op2), .ZN(n1) );
  AND2_X1 U3 ( .A1(op1), .A2(op2), .ZN(g) );
endmodule


module PG_NETWORK_954 ( op1, op2, g, p );
  input op1, op2;
  output g, p;
  wire   n1;

  XNOR2_X1 U1 ( .A(op1), .B(n1), .ZN(p) );
  INV_X1 U2 ( .A(op2), .ZN(n1) );
  AND2_X1 U3 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_953 ( op1, op2, g, p );
  input op1, op2;
  output g, p;
  wire   n1;

  XNOR2_X1 U1 ( .A(n1), .B(op1), .ZN(p) );
  INV_X1 U2 ( .A(op2), .ZN(n1) );
  AND2_X1 U3 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_952 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_951 ( op1, op2, g, p );
  input op1, op2;
  output g, p;
  wire   n1;

  XNOR2_X1 U1 ( .A(op2), .B(n1), .ZN(p) );
  INV_X1 U2 ( .A(op1), .ZN(n1) );
  AND2_X1 U3 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_950 ( op1, op2, g, p );
  input op1, op2;
  output g, p;
  wire   n1;

  AND2_X1 U1 ( .A1(op1), .A2(op2), .ZN(g) );
  XNOR2_X1 U2 ( .A(op2), .B(n1), .ZN(p) );
  INV_X1 U3 ( .A(op1), .ZN(n1) );
endmodule


module PG_NETWORK_949 ( op1, op2, g, p );
  input op1, op2;
  output g, p;
  wire   n1;

  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XNOR2_X1 U2 ( .A(op2), .B(n1), .ZN(p) );
  INV_X1 U3 ( .A(op1), .ZN(n1) );
endmodule


module PG_NETWORK_948 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_947 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op1), .A2(op2), .ZN(g) );
  XOR2_X1 U2 ( .A(op1), .B(op2), .Z(p) );
endmodule


module PG_NETWORK_946 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op1), .B(op2), .Z(p) );
endmodule


module PG_NETWORK_945 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  XOR2_X1 U1 ( .A(op2), .B(op1), .Z(p) );
  AND2_X1 U2 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_944 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_943 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_942 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_941 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  XOR2_X1 U1 ( .A(op1), .B(op2), .Z(p) );
  AND2_X1 U2 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_940 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_939 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_938 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_937 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_936 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_935 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_934 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_933 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_BLOCK_945 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij_BAR );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij_BAR;


  AOI21_X1 U1 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(G_ij_BAR) );
endmodule


module PG_BLOCK_944 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1, n2;

  NAND2_X1 U1 ( .A1(n2), .A2(n1), .ZN(G_ij) );
  INV_X1 U2 ( .A(G_ik), .ZN(n1) );
  NAND2_X1 U3 ( .A1(P_ik), .A2(G_k1j), .ZN(n2) );
  AND2_X1 U4 ( .A1(P_k1j), .A2(P_ik), .ZN(P_ij) );
endmodule


module PG_BLOCK_943 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1, n2;

  NAND2_X1 U1 ( .A1(n2), .A2(n1), .ZN(G_ij) );
  INV_X1 U2 ( .A(G_ik), .ZN(n1) );
  NAND2_X1 U3 ( .A1(P_ik), .A2(G_k1j), .ZN(n2) );
  AND2_X1 U4 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
endmodule


module PG_BLOCK_942 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(G_k1j), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_941 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AOI21_X1 U1 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(G_ij) );
  AND2_X1 U3 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
endmodule


module PG_BLOCK_940 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AOI21_X1 U1 ( .B1(P_ik), .B2(G_k1j), .A(G_ik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(G_ij) );
  AND2_X1 U3 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
endmodule


module PG_BLOCK_939 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1, n2;

  NAND2_X1 U1 ( .A1(n2), .A2(n1), .ZN(G_ij) );
  INV_X1 U2 ( .A(G_ik), .ZN(n1) );
  NAND2_X1 U3 ( .A1(P_ik), .A2(G_k1j), .ZN(n2) );
  AND2_X1 U4 ( .A1(P_k1j), .A2(P_ik), .ZN(P_ij) );
endmodule


module PG_BLOCK_938 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_937 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij_BAR );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij_BAR;


  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(G_ij_BAR) );
endmodule


module PG_BLOCK_936 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_935 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(G_k1j), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_934 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_933 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(G_k1j), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module G_BLOCK_254 ( P_ik, G_k1j, G_ij, G_ik_BAR );
  input P_ik, G_k1j, G_ik_BAR;
  output G_ij;
  wire   G_ik;
  assign G_ik = G_ik_BAR;

  INV_X1 U1 ( .A(G_ik), .ZN(G_ij) );
endmodule


module PG_BLOCK_914 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1, n2;

  NAND2_X1 U1 ( .A1(n2), .A2(n1), .ZN(G_ij) );
  INV_X1 U2 ( .A(G_ik), .ZN(n1) );
  NAND2_X1 U3 ( .A1(P_ik), .A2(G_k1j), .ZN(n2) );
  AND2_X1 U4 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
endmodule


module PG_BLOCK_913 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1, n2;

  NAND2_X1 U1 ( .A1(n2), .A2(n1), .ZN(G_ij) );
  NAND2_X1 U2 ( .A1(G_k1j), .A2(P_ik), .ZN(n1) );
  INV_X1 U3 ( .A(G_ik), .ZN(n2) );
  AND2_X1 U4 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
endmodule


module PG_BLOCK_912 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1, n2;

  NAND2_X1 U1 ( .A1(n2), .A2(n1), .ZN(G_ij) );
  INV_X1 U2 ( .A(G_ik), .ZN(n1) );
  NAND2_X1 U3 ( .A1(G_k1j), .A2(P_ik), .ZN(n2) );
  AND2_X1 U4 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
endmodule


module PG_BLOCK_911 ( P_ik, P_k1j, G_k1j, P_ij, G_ij, G_ik_BAR );
  input P_ik, P_k1j, G_k1j, G_ik_BAR;
  output P_ij, G_ij;
  wire   G_ik, n1;
  assign G_ik = G_ik_BAR;

  NAND2_X1 U1 ( .A1(G_ik), .A2(n1), .ZN(G_ij) );
  NAND2_X1 U2 ( .A1(P_ik), .A2(G_k1j), .ZN(n1) );
  AND2_X1 U3 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
endmodule


module PG_BLOCK_910 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij_BAR );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij_BAR;


  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(G_ij_BAR) );
endmodule


module PG_BLOCK_909 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module G_BLOCK_253 ( P_ik, G_ik, G_k1j, G_ij );
  input P_ik, G_ik, G_k1j;
  output G_ij;
  wire   n1, n2;

  NAND2_X2 U1 ( .A1(n2), .A2(n1), .ZN(G_ij) );
  NAND2_X1 U2 ( .A1(P_ik), .A2(G_k1j), .ZN(n1) );
  INV_X1 U3 ( .A(G_ik), .ZN(n2) );
endmodule


module PG_BLOCK_899 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1, n2;

  NAND2_X1 U1 ( .A1(n2), .A2(n1), .ZN(G_ij) );
  INV_X1 U2 ( .A(G_ik), .ZN(n1) );
  NAND2_X1 U3 ( .A1(G_k1j), .A2(P_ik), .ZN(n2) );
  AND2_X1 U4 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
endmodule


module PG_BLOCK_898 ( P_ik, P_k1j, G_k1j, P_ij, G_ij, G_ik_BAR );
  input P_ik, P_k1j, G_k1j, G_ik_BAR;
  output P_ij, G_ij;
  wire   G_ik, n1;
  assign G_ik = G_ik_BAR;

  NAND2_X1 U1 ( .A1(G_ik), .A2(n1), .ZN(G_ij) );
  NAND2_X1 U2 ( .A1(P_ik), .A2(G_k1j), .ZN(n1) );
  AND2_X1 U3 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
endmodule


module G_BLOCK_252 ( P_ik, G_ik, G_k1j, G_ij );
  input P_ik, G_ik, G_k1j;
  output G_ij;
  wire   n1, n2;

  NAND2_X1 U1 ( .A1(n1), .A2(n2), .ZN(G_ij) );
  NAND2_X1 U2 ( .A1(G_k1j), .A2(P_ik), .ZN(n1) );
  INV_X1 U3 ( .A(G_ik), .ZN(n2) );
endmodule


module G_BLOCK_251 ( P_ik, G_ik, G_k1j, G_ij );
  input P_ik, G_ik, G_k1j;
  output G_ij;
  wire   n1;

  OR2_X2 U1 ( .A1(G_ik), .A2(n1), .ZN(G_ij) );
  AND2_X1 U2 ( .A1(G_k1j), .A2(P_ik), .ZN(n1) );
endmodule


module PG_BLOCK_892 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n2;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n2) );
  INV_X1 U3 ( .A(n2), .ZN(G_ij) );
endmodule


module G_BLOCK_250 ( P_ik, G_ik, G_k1j, G_ij );
  input P_ik, G_ik, G_k1j;
  output G_ij;
  wire   n1, n2;

  NAND2_X1 U1 ( .A1(n2), .A2(n1), .ZN(G_ij) );
  NAND2_X1 U2 ( .A1(G_k1j), .A2(P_ik), .ZN(n1) );
  INV_X1 U3 ( .A(G_ik), .ZN(n2) );
endmodule


module G_BLOCK_249 ( P_ik, G_ik, G_k1j, G_ij );
  input P_ik, G_ik, G_k1j;
  output G_ij;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(G_ij) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(G_k1j), .A(G_ik), .ZN(n2) );
endmodule


module G_BLOCK_248 ( P_ik, G_ik, G_k1j, G_ij );
  input P_ik, G_ik, G_k1j;
  output G_ij;
  wire   n1;

  AOI21_X1 U1 ( .B1(P_ik), .B2(G_k1j), .A(G_ik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(G_ij) );
endmodule


module CARRY_GENERATOR_Nbit64_0 ( A, B, Cin, Cout );
  input [63:0] A;
  input [63:0] B;
  output [16:0] Cout;
  input Cin;
  wire   n8, \p[4][2] , \p[3][2] , \p[3][1] , \p[2][6] , \p[2][5] , \p[2][4] ,
         \p[2][3] , \p[2][2] , \p[2][1] , \p[1][13] , \p[1][12] , \p[1][11] ,
         \p[1][10] , \p[1][9] , \p[1][8] , \p[1][7] , \p[1][6] , \p[1][5] ,
         \p[1][4] , \p[1][3] , \p[1][2] , \p[0][28] , \p[0][27] , \p[0][26] ,
         \p[0][25] , \p[0][24] , \p[0][23] , \p[0][22] , \p[0][21] ,
         \p[0][20] , \p[0][19] , \p[0][18] , \p[0][17] , \p[0][16] ,
         \p[0][15] , \p[0][14] , \p[0][13] , \p[0][12] , \p[0][11] ,
         \p[0][10] , \p[0][9] , \p[0][8] , \p[0][7] , \p[0][6] , \p[0][5] ,
         \p[0][4] , \g[4][2] , \g[3][1] , \g[2][6] , \g[2][5] , \g[2][4] ,
         \g[2][3] , \g[2][2] , \g[2][1] , \g[1][13] , \g[1][12] , \g[1][11] ,
         \g[1][10] , \g[1][9] , \g[1][8] , \g[1][7] , \g[1][6] , \g[1][5] ,
         \g[1][4] , \g[1][3] , \g[1][2] , \g[1][1] , \g[0][28] , \g[0][27] ,
         \g[0][26] , \g[0][25] , \g[0][24] , \g[0][23] , \g[0][22] ,
         \g[0][21] , \g[0][20] , \g[0][19] , \g[0][18] , \g[0][17] ,
         \g[0][16] , \g[0][15] , \g[0][14] , \g[0][13] , \g[0][12] ,
         \g[0][11] , \g[0][10] , \g[0][9] , \g[0][8] , \g[0][7] , \g[0][6] ,
         \g[0][5] , \g[0][4] , \g[0][3] , n2, n3, n4;

  PG_NETWORK_958 Block_PG_NET_3 ( .op1(A[2]), .op2(B[2]), .g(\g[0][3] ) );
  PG_NETWORK_957 Block_PG_NET_4 ( .op1(A[3]), .op2(B[3]), .g(\g[0][4] ), .p(
        \p[0][4] ) );
  PG_NETWORK_956 Block_PG_NET_5 ( .op1(A[4]), .op2(B[4]), .g(\g[0][5] ), .p(
        \p[0][5] ) );
  PG_NETWORK_955 Block_PG_NET_6 ( .op1(A[5]), .op2(B[5]), .g(\g[0][6] ), .p(
        \p[0][6] ) );
  PG_NETWORK_954 Block_PG_NET_7 ( .op1(A[6]), .op2(B[6]), .g(\g[0][7] ), .p(
        \p[0][7] ) );
  PG_NETWORK_953 Block_PG_NET_8 ( .op1(A[7]), .op2(B[7]), .g(\g[0][8] ), .p(
        \p[0][8] ) );
  PG_NETWORK_952 Block_PG_NET_9 ( .op1(A[8]), .op2(B[8]), .g(\g[0][9] ), .p(
        \p[0][9] ) );
  PG_NETWORK_951 Block_PG_NET_10 ( .op1(A[9]), .op2(B[9]), .g(\g[0][10] ), .p(
        \p[0][10] ) );
  PG_NETWORK_950 Block_PG_NET_11 ( .op1(A[10]), .op2(B[10]), .g(\g[0][11] ), 
        .p(\p[0][11] ) );
  PG_NETWORK_949 Block_PG_NET_12 ( .op1(A[11]), .op2(B[11]), .g(\g[0][12] ), 
        .p(\p[0][12] ) );
  PG_NETWORK_948 Block_PG_NET_13 ( .op1(A[12]), .op2(B[12]), .g(\g[0][13] ), 
        .p(\p[0][13] ) );
  PG_NETWORK_947 Block_PG_NET_14 ( .op1(A[13]), .op2(B[13]), .g(\g[0][14] ), 
        .p(\p[0][14] ) );
  PG_NETWORK_946 Block_PG_NET_15 ( .op1(A[14]), .op2(B[14]), .g(\g[0][15] ), 
        .p(\p[0][15] ) );
  PG_NETWORK_945 Block_PG_NET_16 ( .op1(A[15]), .op2(B[15]), .g(\g[0][16] ), 
        .p(\p[0][16] ) );
  PG_NETWORK_944 Block_PG_NET_17 ( .op1(A[16]), .op2(B[16]), .g(\g[0][17] ), 
        .p(\p[0][17] ) );
  PG_NETWORK_943 Block_PG_NET_18 ( .op1(A[17]), .op2(B[17]), .g(\g[0][18] ), 
        .p(\p[0][18] ) );
  PG_NETWORK_942 Block_PG_NET_19 ( .op1(A[18]), .op2(B[18]), .g(\g[0][19] ), 
        .p(\p[0][19] ) );
  PG_NETWORK_941 Block_PG_NET_20 ( .op1(A[19]), .op2(B[19]), .g(\g[0][20] ), 
        .p(\p[0][20] ) );
  PG_NETWORK_940 Block_PG_NET_21 ( .op1(A[20]), .op2(B[20]), .g(\g[0][21] ), 
        .p(\p[0][21] ) );
  PG_NETWORK_939 Block_PG_NET_22 ( .op1(A[21]), .op2(B[21]), .g(\g[0][22] ), 
        .p(\p[0][22] ) );
  PG_NETWORK_938 Block_PG_NET_23 ( .op1(A[22]), .op2(B[22]), .g(\g[0][23] ), 
        .p(\p[0][23] ) );
  PG_NETWORK_937 Block_PG_NET_24 ( .op1(A[23]), .op2(B[23]), .g(\g[0][24] ), 
        .p(\p[0][24] ) );
  PG_NETWORK_936 Block_PG_NET_25 ( .op1(A[24]), .op2(B[24]), .g(\g[0][25] ), 
        .p(\p[0][25] ) );
  PG_NETWORK_935 Block_PG_NET_26 ( .op1(A[25]), .op2(B[25]), .g(\g[0][26] ), 
        .p(\p[0][26] ) );
  PG_NETWORK_934 Block_PG_NET_27 ( .op1(A[26]), .op2(B[26]), .g(\g[0][27] ), 
        .p(\p[0][27] ) );
  PG_NETWORK_933 Block_PG_NET_28 ( .op1(A[27]), .op2(B[27]), .g(\g[0][28] ), 
        .p(\p[0][28] ) );
  PG_BLOCK_945 Block_Stage_ONE_1 ( .P_ik(\p[0][4] ), .G_ik(\g[0][4] ), .P_k1j(
        1'b0), .G_k1j(\g[0][3] ), .G_ij_BAR(\g[1][1] ) );
  PG_BLOCK_944 Block_Stage_ONE_2 ( .P_ik(\p[0][6] ), .G_ik(\g[0][6] ), .P_k1j(
        \p[0][5] ), .G_k1j(\g[0][5] ), .P_ij(\p[1][2] ), .G_ij(\g[1][2] ) );
  PG_BLOCK_943 Block_Stage_ONE_3 ( .P_ik(\p[0][8] ), .G_ik(\g[0][8] ), .P_k1j(
        \p[0][7] ), .G_k1j(\g[0][7] ), .P_ij(\p[1][3] ), .G_ij(\g[1][3] ) );
  PG_BLOCK_942 Block_Stage_ONE_4 ( .P_ik(\p[0][10] ), .G_ik(\g[0][10] ), 
        .P_k1j(\p[0][9] ), .G_k1j(\g[0][9] ), .P_ij(\p[1][4] ), .G_ij(
        \g[1][4] ) );
  PG_BLOCK_941 Block_Stage_ONE_5 ( .P_ik(\p[0][12] ), .G_ik(\g[0][12] ), 
        .P_k1j(\p[0][11] ), .G_k1j(\g[0][11] ), .P_ij(\p[1][5] ), .G_ij(
        \g[1][5] ) );
  PG_BLOCK_940 Block_Stage_ONE_6 ( .P_ik(\p[0][14] ), .G_ik(\g[0][14] ), 
        .P_k1j(\p[0][13] ), .G_k1j(\g[0][13] ), .P_ij(\p[1][6] ), .G_ij(
        \g[1][6] ) );
  PG_BLOCK_939 Block_Stage_ONE_7 ( .P_ik(\p[0][16] ), .G_ik(\g[0][16] ), 
        .P_k1j(\p[0][15] ), .G_k1j(\g[0][15] ), .P_ij(\p[1][7] ), .G_ij(
        \g[1][7] ) );
  PG_BLOCK_938 Block_Stage_ONE_8 ( .P_ik(\p[0][18] ), .G_ik(\g[0][18] ), 
        .P_k1j(\p[0][17] ), .G_k1j(\g[0][17] ), .P_ij(\p[1][8] ), .G_ij(
        \g[1][8] ) );
  PG_BLOCK_937 Block_Stage_ONE_9 ( .P_ik(\p[0][20] ), .G_ik(\g[0][20] ), 
        .P_k1j(\p[0][19] ), .G_k1j(\g[0][19] ), .P_ij(\p[1][9] ), .G_ij_BAR(
        \g[1][9] ) );
  PG_BLOCK_936 Block_Stage_ONE_10 ( .P_ik(\p[0][22] ), .G_ik(\g[0][22] ), 
        .P_k1j(\p[0][21] ), .G_k1j(\g[0][21] ), .P_ij(\p[1][10] ), .G_ij(
        \g[1][10] ) );
  PG_BLOCK_935 Block_Stage_ONE_11 ( .P_ik(\p[0][24] ), .G_ik(\g[0][24] ), 
        .P_k1j(\p[0][23] ), .G_k1j(\g[0][23] ), .P_ij(\p[1][11] ), .G_ij(
        \g[1][11] ) );
  PG_BLOCK_934 Block_Stage_ONE_12 ( .P_ik(\p[0][26] ), .G_ik(\g[0][26] ), 
        .P_k1j(\p[0][25] ), .G_k1j(\g[0][25] ), .P_ij(\p[1][12] ), .G_ij(
        \g[1][12] ) );
  PG_BLOCK_933 Block_Stage_ONE_13 ( .P_ik(\p[0][28] ), .G_ik(\g[0][28] ), 
        .P_k1j(\p[0][27] ), .G_k1j(\g[0][27] ), .P_ij(\p[1][13] ), .G_ij(
        \g[1][13] ) );
  G_BLOCK_254 g_2 ( .P_ik(1'b0), .G_k1j(1'b0), .G_ij(n8), .G_ik_BAR(\g[1][1] )
         );
  PG_BLOCK_914 Block_Stage_TWO_1 ( .P_ik(\p[1][3] ), .G_ik(\g[1][3] ), .P_k1j(
        \p[1][2] ), .G_k1j(\g[1][2] ), .P_ij(\p[2][1] ), .G_ij(\g[2][1] ) );
  PG_BLOCK_913 Block_Stage_TWO_2 ( .P_ik(\p[1][5] ), .G_ik(\g[1][5] ), .P_k1j(
        \p[1][4] ), .G_k1j(\g[1][4] ), .P_ij(\p[2][2] ), .G_ij(\g[2][2] ) );
  PG_BLOCK_912 Block_Stage_TWO_3 ( .P_ik(\p[1][7] ), .G_ik(\g[1][7] ), .P_k1j(
        \p[1][6] ), .G_k1j(\g[1][6] ), .P_ij(\p[2][3] ), .G_ij(\g[2][3] ) );
  PG_BLOCK_911 Block_Stage_TWO_4 ( .P_ik(\p[1][9] ), .P_k1j(\p[1][8] ), 
        .G_k1j(\g[1][8] ), .P_ij(\p[2][4] ), .G_ij(\g[2][4] ), .G_ik_BAR(
        \g[1][9] ) );
  PG_BLOCK_910 Block_Stage_TWO_5 ( .P_ik(\p[1][11] ), .G_ik(\g[1][11] ), 
        .P_k1j(\p[1][10] ), .G_k1j(\g[1][10] ), .P_ij(\p[2][5] ), .G_ij_BAR(
        \g[2][5] ) );
  PG_BLOCK_909 Block_Stage_TWO_6 ( .P_ik(\p[1][13] ), .G_ik(\g[1][13] ), 
        .P_k1j(\p[1][12] ), .G_k1j(\g[1][12] ), .P_ij(\p[2][6] ), .G_ij(
        \g[2][6] ) );
  G_BLOCK_253 g_3 ( .P_ik(\p[2][1] ), .G_ik(\g[2][1] ), .G_k1j(n8), .G_ij(
        Cout[2]) );
  PG_BLOCK_899 Block_Stage_THREE_1 ( .P_ik(\p[2][3] ), .G_ik(\g[2][3] ), 
        .P_k1j(\p[2][2] ), .G_k1j(\g[2][2] ), .P_ij(\p[3][1] ), .G_ij(
        \g[3][1] ) );
  PG_BLOCK_898 Block_Stage_THREE_2 ( .P_ik(\p[2][5] ), .P_k1j(\p[2][4] ), 
        .G_k1j(\g[2][4] ), .P_ij(\p[3][2] ), .G_ij(n2), .G_ik_BAR(\g[2][5] )
         );
  G_BLOCK_252 g_4_c12_c16_0 ( .P_ik(\p[2][2] ), .G_ik(\g[2][2] ), .G_k1j(
        Cout[2]), .G_ij(Cout[3]) );
  G_BLOCK_251 g_4_c12_c16_1 ( .P_ik(\p[3][1] ), .G_ik(\g[3][1] ), .G_k1j(
        Cout[2]), .G_ij(Cout[4]) );
  PG_BLOCK_892 Block_stage_FOUR_2_0 ( .P_ik(\p[2][6] ), .G_ik(\g[2][6] ), 
        .P_k1j(\p[3][2] ), .G_k1j(n2), .P_ij(\p[4][2] ), .G_ij(\g[4][2] ) );
  G_BLOCK_250 Block_stage_FIVE_4 ( .P_ik(\p[2][4] ), .G_ik(\g[2][4] ), .G_k1j(
        Cout[4]), .G_ij(Cout[5]) );
  G_BLOCK_249 Block_stage_FIVE_5 ( .P_ik(\p[3][2] ), .G_ik(n2), .G_k1j(n4), 
        .G_ij(Cout[6]) );
  G_BLOCK_248 Block_stage_FIVE_6 ( .P_ik(\p[4][2] ), .G_ik(\g[4][2] ), .G_k1j(
        n4), .G_ij(Cout[7]) );
  BUF_X1 U1 ( .A(n8), .Z(Cout[1]) );
  INV_X1 U2 ( .A(Cout[4]), .ZN(n3) );
  INV_X1 U3 ( .A(n3), .ZN(n4) );
endmodule


module FA_1920 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1919 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1918 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1917 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_480 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \CTMP[3] ;

  FA_1920 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_1919 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_1918 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(1'b0), .S(S[2]), .Co(\CTMP[3] ) );
  FA_1917 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(\CTMP[3] ), .S(S[3]) );
endmodule


module MUX_2to1_N4_240 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_240 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_480 RCA_0 ( .A({A[3:2], 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0) );
  MUX_2to1_N4_240 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_1912 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1911 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(B), .B(A), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1910 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1909 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_478 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1912 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1911 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1910 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1909 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1908 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_1907 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(B), .B(A), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1906 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1905 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_477 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1908 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1907 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1906 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1905 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_239 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;
  wire   n1, n2, n3;

  INV_X1 U1 ( .A(SEL), .ZN(n2) );
  NAND2_X1 U2 ( .A1(n3), .A2(n1), .ZN(Y[3]) );
  NAND2_X1 U3 ( .A1(IN0[3]), .A2(n2), .ZN(n1) );
  NAND2_X1 U4 ( .A1(IN1[3]), .A2(SEL), .ZN(n3) );
  MUX2_X1 U5 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U6 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U7 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
endmodule


module carry_select_block_N4_239 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_478 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_477 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_239 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_1904 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  BUF_X1 U1 ( .A(B), .Z(n1) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U3 ( .A(n1), .B(A), .Z(S) );
endmodule


module FA_1903 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1902 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1901 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(Ci), .B(n1), .ZN(S) );
endmodule


module RCA_N4_476 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1904 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1903 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1902 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1901 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1900 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_1899 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4;

  OR2_X1 U1 ( .A1(B), .A2(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(B), .B(Ci), .ZN(n1) );
  XNOR2_X1 U3 ( .A(n1), .B(A), .ZN(S) );
  NAND2_X1 U4 ( .A1(n3), .A2(n2), .ZN(Co) );
  NAND2_X1 U5 ( .A1(B), .A2(A), .ZN(n2) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n4), .ZN(n3) );
endmodule


module FA_1898 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n1) );
  XOR2_X1 U2 ( .A(Ci), .B(n1), .Z(S) );
  NAND2_X1 U3 ( .A1(Ci), .A2(B), .ZN(n2) );
  NAND2_X1 U4 ( .A1(Ci), .A2(A), .ZN(n3) );
  NAND2_X1 U5 ( .A1(B), .A2(A), .ZN(n4) );
  NAND3_X1 U6 ( .A1(n2), .A2(n3), .A3(n4), .ZN(Co) );
endmodule


module FA_1897 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_475 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1900 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1899 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1898 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1897 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_238 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X2 U2 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
  MUX2_X1 U3 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U4 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
endmodule


module carry_select_block_N4_238 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_476 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_475 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_238 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_1896 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1895 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1894 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1893 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_474 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1896 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1895 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1894 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1893 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1892 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_1891 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1890 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3;

  XNOR2_X1 U1 ( .A(Ci), .B(A), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(B), .ZN(S) );
  INV_X1 U3 ( .A(n2), .ZN(Co) );
  AOI22_X1 U4 ( .A1(Ci), .A2(n3), .B1(B), .B2(A), .ZN(n2) );
  OR2_X1 U5 ( .A1(A), .A2(B), .ZN(n3) );
endmodule


module FA_1889 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_473 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1892 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1891 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1890 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1889 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_237 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U2 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U3 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U4 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
endmodule


module carry_select_block_N4_237 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_474 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_473 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_237 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_1888 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1887 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1886 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1885 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_472 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1888 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1887 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1886 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1885 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1884 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_1883 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(Ci), .CI(B), .CO(Co), .S(S) );
endmodule


module FA_1882 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1881 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_471 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1884 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1883 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1882 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1881 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_236 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
  MUX2_X1 U2 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U3 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U4 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
endmodule


module carry_select_block_N4_236 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_472 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_471 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_236 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_1880 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1879 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1878 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1877 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_470 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1880 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1879 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1878 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1877 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1876 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(S) );
endmodule


module FA_1875 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1874 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1873 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(Ci), .B(n1), .ZN(S) );
endmodule


module RCA_N4_469 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1876 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1875 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1874 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1873 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_235 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
  MUX2_X1 U2 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U3 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U4 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
endmodule


module carry_select_block_N4_235 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_470 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_469 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_235 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_1872 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(S) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(Co) );
endmodule


module FA_1871 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1870 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1869 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(Ci), .B(n1), .ZN(S) );
endmodule


module RCA_N4_468 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1872 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1871 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1870 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1869 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1868 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(S) );
  OR2_X1 U2 ( .A1(A), .A2(B), .ZN(Co) );
endmodule


module FA_1867 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1866 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3;

  OAI21_X1 U1 ( .B1(A), .B2(B), .A(Ci), .ZN(n3) );
  XNOR2_X1 U2 ( .A(Ci), .B(n1), .ZN(S) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n1) );
  NAND2_X1 U4 ( .A1(n3), .A2(n2), .ZN(Co) );
  NAND2_X1 U5 ( .A1(B), .A2(A), .ZN(n2) );
endmodule


module FA_1865 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(Ci), .B(n1), .ZN(S) );
endmodule


module RCA_N4_467 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1868 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1867 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1866 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1865 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_234 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
  MUX2_X1 U3 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X2 U4 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
endmodule


module carry_select_block_N4_234 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_468 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_467 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_234 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_1864 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(S) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(Co) );
endmodule


module FA_1863 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1862 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1861 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_466 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1864 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1863 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1862 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1861 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1860 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(S) );
  OR2_X1 U2 ( .A1(A), .A2(B), .ZN(Co) );
endmodule


module FA_1859 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1858 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1857 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_465 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1860 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1859 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1858 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1857 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_233 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U3 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U4 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
endmodule


module carry_select_block_N4_233 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_466 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_465 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_233 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module SUMGENERATOR_Nblocks16_bits_per_block4_0 ( A, B, CARRY_SELECT, SUM );
  input [63:0] A;
  input [63:0] B;
  input [15:0] CARRY_SELECT;
  output [63:0] SUM;


  carry_select_block_N4_240 block_n_1 ( .A({A[3:2], 1'b0, 1'b0}), .B(B[3:0]), 
        .S(SUM[3:0]), .Ci(1'b0) );
  carry_select_block_N4_239 block_n_2 ( .A(A[7:4]), .B(B[7:4]), .S(SUM[7:4]), 
        .Ci(CARRY_SELECT[1]) );
  carry_select_block_N4_238 block_n_3 ( .A(A[11:8]), .B(B[11:8]), .S(SUM[11:8]), .Ci(CARRY_SELECT[2]) );
  carry_select_block_N4_237 block_n_4 ( .A(A[15:12]), .B(B[15:12]), .S(
        SUM[15:12]), .Ci(CARRY_SELECT[3]) );
  carry_select_block_N4_236 block_n_5 ( .A(A[19:16]), .B(B[19:16]), .S(
        SUM[19:16]), .Ci(CARRY_SELECT[4]) );
  carry_select_block_N4_235 block_n_6 ( .A(A[23:20]), .B(B[23:20]), .S(
        SUM[23:20]), .Ci(CARRY_SELECT[5]) );
  carry_select_block_N4_234 block_n_7 ( .A(A[27:24]), .B(B[27:24]), .S(
        SUM[27:24]), .Ci(CARRY_SELECT[6]) );
  carry_select_block_N4_233 block_n_8 ( .A(A[31:28]), .B(B[31:28]), .S(
        SUM[31:28]), .Ci(CARRY_SELECT[7]) );
endmodule


module ADDER_P4_N_BIT64_0 ( A, B, add_sub, Cout, SUM );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input add_sub;
  output Cout;
  wire   n1, n2, n3;
  wire   [63:0] B_xor;
  wire   [15:0] tmp_co;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41;
  assign B_xor[31] = B[31];
  assign B_xor[30] = B[30];
  assign B_xor[29] = B[29];
  assign B_xor[28] = B[28];
  assign B_xor[27] = B[27];
  assign B_xor[26] = B[26];
  assign B_xor[25] = B[25];
  assign B_xor[24] = B[24];
  assign B_xor[23] = B[23];
  assign B_xor[22] = B[22];
  assign B_xor[21] = B[21];
  assign B_xor[20] = B[20];
  assign B_xor[19] = B[19];
  assign B_xor[18] = B[18];
  assign B_xor[17] = B[17];
  assign B_xor[16] = B[16];
  assign B_xor[15] = B[15];
  assign B_xor[14] = B[14];
  assign B_xor[13] = B[13];
  assign B_xor[12] = B[12];
  assign B_xor[11] = B[11];
  assign B_xor[10] = B[10];
  assign B_xor[9] = B[9];
  assign B_xor[8] = B[8];
  assign B_xor[7] = B[7];
  assign B_xor[6] = B[6];
  assign B_xor[5] = B[5];
  assign B_xor[4] = B[4];
  assign B_xor[3] = B[3];
  assign B_xor[2] = B[2];
  assign B_xor[1] = B[1];
  assign B_xor[0] = B[0];

  CARRY_GENERATOR_Nbit64_0 CLA_SPARSE_TREE ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, A[27:2], 1'b0, 1'b0}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        B_xor[27:2], 1'b0, 1'b0}), .Cin(1'b0), .Cout({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, tmp_co[7:1], 
        SYNOPSYS_UNCONNECTED__9}) );
  SUMGENERATOR_Nblocks16_bits_per_block4_0 CSA ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, A[31:8], n1, A[6], n3, A[4:2], 1'b0, 1'b0}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B_xor[31:0]}), 
        .CARRY_SELECT({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        tmp_co[7:1], 1'b0}), .SUM({SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, SYNOPSYS_UNCONNECTED__22, 
        SYNOPSYS_UNCONNECTED__23, SYNOPSYS_UNCONNECTED__24, 
        SYNOPSYS_UNCONNECTED__25, SYNOPSYS_UNCONNECTED__26, 
        SYNOPSYS_UNCONNECTED__27, SYNOPSYS_UNCONNECTED__28, 
        SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, 
        SYNOPSYS_UNCONNECTED__31, SYNOPSYS_UNCONNECTED__32, 
        SYNOPSYS_UNCONNECTED__33, SYNOPSYS_UNCONNECTED__34, 
        SYNOPSYS_UNCONNECTED__35, SYNOPSYS_UNCONNECTED__36, 
        SYNOPSYS_UNCONNECTED__37, SYNOPSYS_UNCONNECTED__38, 
        SYNOPSYS_UNCONNECTED__39, SYNOPSYS_UNCONNECTED__40, 
        SYNOPSYS_UNCONNECTED__41, SUM[31:0]}) );
  BUF_X1 U1 ( .A(A[7]), .Z(n1) );
  INV_X1 U2 ( .A(A[5]), .ZN(n2) );
  INV_X1 U3 ( .A(n2), .ZN(n3) );
endmodule


module PG_NETWORK_892 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_891 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_890 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_889 ( op1, op2, g, p );
  input op1, op2;
  output g, p;
  wire   n1;

  XNOR2_X1 U1 ( .A(op2), .B(n1), .ZN(p) );
  INV_X1 U2 ( .A(op1), .ZN(n1) );
  AND2_X1 U3 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_888 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_887 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_886 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_885 ( op1, op2, g, p );
  input op1, op2;
  output g, p;
  wire   n1;

  XNOR2_X1 U1 ( .A(op2), .B(n1), .ZN(p) );
  INV_X1 U2 ( .A(op1), .ZN(n1) );
  AND2_X1 U3 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_884 ( op1, op2, g, p );
  input op1, op2;
  output g, p;
  wire   n1;

  XNOR2_X1 U1 ( .A(op2), .B(n1), .ZN(p) );
  INV_X1 U2 ( .A(op1), .ZN(n1) );
  AND2_X1 U3 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_883 ( op1, op2, g, p );
  input op1, op2;
  output g, p;
  wire   n1;

  XNOR2_X1 U1 ( .A(op2), .B(n1), .ZN(p) );
  INV_X1 U2 ( .A(op1), .ZN(n1) );
  AND2_X1 U3 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_882 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_881 ( op1, op2, g, p );
  input op1, op2;
  output g, p;
  wire   n1;

  XNOR2_X1 U1 ( .A(op2), .B(n1), .ZN(p) );
  INV_X1 U2 ( .A(op1), .ZN(n1) );
  AND2_X1 U3 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_880 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_879 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_878 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_877 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_876 ( op1, op2, g, p );
  input op1, op2;
  output g, p;
  wire   n1;

  XNOR2_X1 U1 ( .A(op2), .B(n1), .ZN(p) );
  INV_X1 U2 ( .A(op1), .ZN(n1) );
  AND2_X1 U3 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_875 ( op1, op2, g, p );
  input op1, op2;
  output g, p;
  wire   n1;

  XNOR2_X1 U1 ( .A(op2), .B(n1), .ZN(p) );
  INV_X1 U2 ( .A(op1), .ZN(n1) );
  AND2_X1 U3 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_874 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_873 ( op1, op2, g, p );
  input op1, op2;
  output g, p;
  wire   n1;

  XNOR2_X1 U1 ( .A(op2), .B(n1), .ZN(p) );
  INV_X1 U2 ( .A(op1), .ZN(n1) );
  AND2_X1 U3 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_872 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_871 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_870 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_869 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_BLOCK_881 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AOI21_X1 U1 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_880 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(G_k1j), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_879 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_878 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1, n2;

  NAND2_X1 U1 ( .A1(n2), .A2(n1), .ZN(G_ij) );
  INV_X1 U2 ( .A(G_ik), .ZN(n1) );
  NAND2_X1 U3 ( .A1(P_ik), .A2(G_k1j), .ZN(n2) );
  AND2_X1 U4 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
endmodule


module PG_BLOCK_877 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1, n2;

  NAND2_X1 U1 ( .A1(n2), .A2(n1), .ZN(G_ij) );
  INV_X1 U2 ( .A(G_ik), .ZN(n1) );
  NAND2_X1 U3 ( .A1(P_ik), .A2(G_k1j), .ZN(n2) );
  AND2_X1 U4 ( .A1(P_k1j), .A2(P_ik), .ZN(P_ij) );
endmodule


module PG_BLOCK_876 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1, n2;

  NAND2_X1 U1 ( .A1(n2), .A2(n1), .ZN(G_ij) );
  INV_X1 U2 ( .A(G_ik), .ZN(n1) );
  NAND2_X1 U3 ( .A1(P_ik), .A2(G_k1j), .ZN(n2) );
  AND2_X1 U4 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
endmodule


module PG_BLOCK_875 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_874 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(G_k1j), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_873 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1, n2;

  NAND2_X1 U1 ( .A1(n2), .A2(n1), .ZN(G_ij) );
  INV_X1 U2 ( .A(G_ik), .ZN(n1) );
  NAND2_X1 U3 ( .A1(P_ik), .A2(G_k1j), .ZN(n2) );
  AND2_X1 U4 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
endmodule


module PG_BLOCK_872 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1, n2;

  NAND2_X1 U1 ( .A1(n2), .A2(n1), .ZN(G_ij) );
  INV_X1 U2 ( .A(G_ik), .ZN(n1) );
  NAND2_X1 U3 ( .A1(P_ik), .A2(G_k1j), .ZN(n2) );
  AND2_X1 U4 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
endmodule


module PG_BLOCK_871 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_k1j), .A2(P_ik), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_870 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij_BAR );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij_BAR;


  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(G_k1j), .A(G_ik), .ZN(G_ij_BAR) );
endmodule


module PG_BLOCK_851 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij_BAR );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij_BAR;
  wire   n1;

  NOR2_X1 U1 ( .A1(n1), .A2(G_ik), .ZN(G_ij_BAR) );
  AND2_X1 U2 ( .A1(P_ik), .A2(G_k1j), .ZN(n1) );
endmodule


module PG_BLOCK_850 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_849 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1, n2;

  NAND2_X1 U1 ( .A1(n2), .A2(n1), .ZN(G_ij) );
  INV_X1 U2 ( .A(G_ik), .ZN(n1) );
  NAND2_X1 U3 ( .A1(G_k1j), .A2(P_ik), .ZN(n2) );
  AND2_X1 U4 ( .A1(P_k1j), .A2(P_ik), .ZN(P_ij) );
endmodule


module PG_BLOCK_848 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_847 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1, n2;

  NAND2_X1 U1 ( .A1(n1), .A2(n2), .ZN(G_ij) );
  INV_X1 U2 ( .A(G_ik), .ZN(n1) );
  NAND2_X1 U3 ( .A1(G_k1j), .A2(P_ik), .ZN(n2) );
  AND2_X1 U4 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
endmodule


module PG_BLOCK_846 ( P_ik, P_k1j, G_k1j, P_ij, G_ij, G_ik_BAR );
  input P_ik, P_k1j, G_k1j, G_ik_BAR;
  output P_ij, G_ij;
  wire   G_ik, n1;
  assign G_ik = G_ik_BAR;

  NAND2_X1 U1 ( .A1(n1), .A2(G_ik), .ZN(G_ij) );
  NAND2_X1 U2 ( .A1(G_k1j), .A2(P_ik), .ZN(n1) );
  AND2_X1 U3 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
endmodule


module G_BLOCK_236 ( P_ik, G_k1j, G_ij, G_ik_BAR );
  input P_ik, G_k1j, G_ik_BAR;
  output G_ij;
  wire   G_ik;
  assign G_ik = G_ik_BAR;

  INV_X1 U1 ( .A(G_ik), .ZN(G_ij) );
endmodule


module PG_BLOCK_836 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1, n2;

  NAND2_X1 U1 ( .A1(n2), .A2(n1), .ZN(G_ij) );
  NAND2_X1 U2 ( .A1(P_ik), .A2(G_k1j), .ZN(n1) );
  INV_X1 U3 ( .A(G_ik), .ZN(n2) );
  AND2_X1 U4 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
endmodule


module PG_BLOCK_835 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1, n2;

  NAND2_X1 U1 ( .A1(n2), .A2(n1), .ZN(G_ij) );
  NAND2_X1 U2 ( .A1(P_ik), .A2(G_k1j), .ZN(n1) );
  INV_X1 U3 ( .A(G_ik), .ZN(n2) );
  AND2_X1 U4 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
endmodule


module G_BLOCK_235 ( P_ik, G_ik, G_k1j, G_ij );
  input P_ik, G_ik, G_k1j;
  output G_ij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(G_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
endmodule


module G_BLOCK_234 ( P_ik, G_ik, G_k1j, G_ij );
  input P_ik, G_ik, G_k1j;
  output G_ij;
  wire   n1;

  OR2_X2 U1 ( .A1(n1), .A2(G_ik), .ZN(G_ij) );
  AND2_X1 U2 ( .A1(P_ik), .A2(G_k1j), .ZN(n1) );
endmodule


module PG_BLOCK_829 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1, n2;

  NAND2_X1 U1 ( .A1(n2), .A2(n1), .ZN(G_ij) );
  NAND2_X1 U2 ( .A1(P_ik), .A2(G_k1j), .ZN(n1) );
  INV_X1 U3 ( .A(G_ik), .ZN(n2) );
  AND2_X1 U4 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
endmodule


module G_BLOCK_233 ( P_ik, G_ik, G_k1j, G_ij );
  input P_ik, G_ik, G_k1j;
  output G_ij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(G_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
endmodule


module G_BLOCK_232 ( P_ik, G_ik, G_k1j, G_ij );
  input P_ik, G_ik, G_k1j;
  output G_ij;
  wire   n1;

  OR2_X2 U1 ( .A1(G_ik), .A2(n1), .ZN(G_ij) );
  AND2_X1 U2 ( .A1(G_k1j), .A2(P_ik), .ZN(n1) );
endmodule


module G_BLOCK_231 ( P_ik, G_ik, G_k1j, G_ij );
  input P_ik, G_ik, G_k1j;
  output G_ij;
  wire   n1;

  AOI21_X1 U1 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(G_ij) );
endmodule


module CARRY_GENERATOR_Nbit64_14 ( A, B, Cin, Cout );
  input [63:0] A;
  input [63:0] B;
  output [16:0] Cout;
  input Cin;
  wire   \p[4][2] , \p[3][2] , \p[3][1] , \p[2][6] , \p[2][5] , \p[2][4] ,
         \p[2][3] , \p[2][2] , \p[1][13] , \p[1][12] , \p[1][11] , \p[1][10] ,
         \p[1][9] , \p[1][8] , \p[1][7] , \p[1][6] , \p[1][5] , \p[1][4] ,
         \p[1][3] , \p[0][28] , \p[0][27] , \p[0][26] , \p[0][25] , \p[0][24] ,
         \p[0][23] , \p[0][22] , \p[0][21] , \p[0][20] , \p[0][19] ,
         \p[0][18] , \p[0][17] , \p[0][16] , \p[0][15] , \p[0][14] ,
         \p[0][13] , \p[0][12] , \p[0][11] , \p[0][10] , \p[0][9] , \p[0][8] ,
         \p[0][7] , \p[0][6] , \g[4][2] , \g[3][2] , \g[3][1] , \g[2][6] ,
         \g[2][5] , \g[2][4] , \g[2][3] , \g[2][2] , \g[2][1] , \g[1][13] ,
         \g[1][12] , \g[1][11] , \g[1][10] , \g[1][9] , \g[1][8] , \g[1][7] ,
         \g[1][6] , \g[1][5] , \g[1][4] , \g[1][3] , \g[1][2] , \g[0][28] ,
         \g[0][27] , \g[0][26] , \g[0][25] , \g[0][24] , \g[0][23] ,
         \g[0][22] , \g[0][21] , \g[0][20] , \g[0][19] , \g[0][18] ,
         \g[0][17] , \g[0][16] , \g[0][15] , \g[0][14] , \g[0][13] ,
         \g[0][12] , \g[0][11] , \g[0][10] , \g[0][9] , \g[0][8] , \g[0][7] ,
         \g[0][6] , \g[0][5] ;

  PG_NETWORK_892 Block_PG_NET_5 ( .op1(A[4]), .op2(B[4]), .g(\g[0][5] ) );
  PG_NETWORK_891 Block_PG_NET_6 ( .op1(A[5]), .op2(B[5]), .g(\g[0][6] ), .p(
        \p[0][6] ) );
  PG_NETWORK_890 Block_PG_NET_7 ( .op1(A[6]), .op2(B[6]), .g(\g[0][7] ), .p(
        \p[0][7] ) );
  PG_NETWORK_889 Block_PG_NET_8 ( .op1(A[7]), .op2(B[7]), .g(\g[0][8] ), .p(
        \p[0][8] ) );
  PG_NETWORK_888 Block_PG_NET_9 ( .op1(A[8]), .op2(B[8]), .g(\g[0][9] ), .p(
        \p[0][9] ) );
  PG_NETWORK_887 Block_PG_NET_10 ( .op1(A[9]), .op2(B[9]), .g(\g[0][10] ), .p(
        \p[0][10] ) );
  PG_NETWORK_886 Block_PG_NET_11 ( .op1(A[10]), .op2(B[10]), .g(\g[0][11] ), 
        .p(\p[0][11] ) );
  PG_NETWORK_885 Block_PG_NET_12 ( .op1(A[11]), .op2(B[11]), .g(\g[0][12] ), 
        .p(\p[0][12] ) );
  PG_NETWORK_884 Block_PG_NET_13 ( .op1(A[12]), .op2(B[12]), .g(\g[0][13] ), 
        .p(\p[0][13] ) );
  PG_NETWORK_883 Block_PG_NET_14 ( .op1(A[13]), .op2(B[13]), .g(\g[0][14] ), 
        .p(\p[0][14] ) );
  PG_NETWORK_882 Block_PG_NET_15 ( .op1(A[14]), .op2(B[14]), .g(\g[0][15] ), 
        .p(\p[0][15] ) );
  PG_NETWORK_881 Block_PG_NET_16 ( .op1(A[15]), .op2(B[15]), .g(\g[0][16] ), 
        .p(\p[0][16] ) );
  PG_NETWORK_880 Block_PG_NET_17 ( .op1(A[16]), .op2(B[16]), .g(\g[0][17] ), 
        .p(\p[0][17] ) );
  PG_NETWORK_879 Block_PG_NET_18 ( .op1(A[17]), .op2(B[17]), .g(\g[0][18] ), 
        .p(\p[0][18] ) );
  PG_NETWORK_878 Block_PG_NET_19 ( .op1(A[18]), .op2(B[18]), .g(\g[0][19] ), 
        .p(\p[0][19] ) );
  PG_NETWORK_877 Block_PG_NET_20 ( .op1(A[19]), .op2(B[19]), .g(\g[0][20] ), 
        .p(\p[0][20] ) );
  PG_NETWORK_876 Block_PG_NET_21 ( .op1(A[20]), .op2(B[20]), .g(\g[0][21] ), 
        .p(\p[0][21] ) );
  PG_NETWORK_875 Block_PG_NET_22 ( .op1(A[21]), .op2(B[21]), .g(\g[0][22] ), 
        .p(\p[0][22] ) );
  PG_NETWORK_874 Block_PG_NET_23 ( .op1(A[22]), .op2(B[22]), .g(\g[0][23] ), 
        .p(\p[0][23] ) );
  PG_NETWORK_873 Block_PG_NET_24 ( .op1(A[23]), .op2(B[23]), .g(\g[0][24] ), 
        .p(\p[0][24] ) );
  PG_NETWORK_872 Block_PG_NET_25 ( .op1(A[24]), .op2(B[24]), .g(\g[0][25] ), 
        .p(\p[0][25] ) );
  PG_NETWORK_871 Block_PG_NET_26 ( .op1(A[25]), .op2(B[25]), .g(\g[0][26] ), 
        .p(\p[0][26] ) );
  PG_NETWORK_870 Block_PG_NET_27 ( .op1(A[26]), .op2(B[26]), .g(\g[0][27] ), 
        .p(\p[0][27] ) );
  PG_NETWORK_869 Block_PG_NET_28 ( .op1(A[27]), .op2(B[27]), .g(\g[0][28] ), 
        .p(\p[0][28] ) );
  PG_BLOCK_881 Block_Stage_ONE_2 ( .P_ik(\p[0][6] ), .G_ik(\g[0][6] ), .P_k1j(
        1'b0), .G_k1j(\g[0][5] ), .G_ij(\g[1][2] ) );
  PG_BLOCK_880 Block_Stage_ONE_3 ( .P_ik(\p[0][8] ), .G_ik(\g[0][8] ), .P_k1j(
        \p[0][7] ), .G_k1j(\g[0][7] ), .P_ij(\p[1][3] ), .G_ij(\g[1][3] ) );
  PG_BLOCK_879 Block_Stage_ONE_4 ( .P_ik(\p[0][10] ), .G_ik(\g[0][10] ), 
        .P_k1j(\p[0][9] ), .G_k1j(\g[0][9] ), .P_ij(\p[1][4] ), .G_ij(
        \g[1][4] ) );
  PG_BLOCK_878 Block_Stage_ONE_5 ( .P_ik(\p[0][12] ), .G_ik(\g[0][12] ), 
        .P_k1j(\p[0][11] ), .G_k1j(\g[0][11] ), .P_ij(\p[1][5] ), .G_ij(
        \g[1][5] ) );
  PG_BLOCK_877 Block_Stage_ONE_6 ( .P_ik(\p[0][14] ), .G_ik(\g[0][14] ), 
        .P_k1j(\p[0][13] ), .G_k1j(\g[0][13] ), .P_ij(\p[1][6] ), .G_ij(
        \g[1][6] ) );
  PG_BLOCK_876 Block_Stage_ONE_7 ( .P_ik(\p[0][16] ), .G_ik(\g[0][16] ), 
        .P_k1j(\p[0][15] ), .G_k1j(\g[0][15] ), .P_ij(\p[1][7] ), .G_ij(
        \g[1][7] ) );
  PG_BLOCK_875 Block_Stage_ONE_8 ( .P_ik(\p[0][18] ), .G_ik(\g[0][18] ), 
        .P_k1j(\p[0][17] ), .G_k1j(\g[0][17] ), .P_ij(\p[1][8] ), .G_ij(
        \g[1][8] ) );
  PG_BLOCK_874 Block_Stage_ONE_9 ( .P_ik(\p[0][20] ), .G_ik(\g[0][20] ), 
        .P_k1j(\p[0][19] ), .G_k1j(\g[0][19] ), .P_ij(\p[1][9] ), .G_ij(
        \g[1][9] ) );
  PG_BLOCK_873 Block_Stage_ONE_10 ( .P_ik(\p[0][22] ), .G_ik(\g[0][22] ), 
        .P_k1j(\p[0][21] ), .G_k1j(\g[0][21] ), .P_ij(\p[1][10] ), .G_ij(
        \g[1][10] ) );
  PG_BLOCK_872 Block_Stage_ONE_11 ( .P_ik(\p[0][24] ), .G_ik(\g[0][24] ), 
        .P_k1j(\p[0][23] ), .G_k1j(\g[0][23] ), .P_ij(\p[1][11] ), .G_ij(
        \g[1][11] ) );
  PG_BLOCK_871 Block_Stage_ONE_12 ( .P_ik(\p[0][26] ), .G_ik(\g[0][26] ), 
        .P_k1j(\p[0][25] ), .G_k1j(\g[0][25] ), .P_ij(\p[1][12] ), .G_ij(
        \g[1][12] ) );
  PG_BLOCK_870 Block_Stage_ONE_13 ( .P_ik(\p[0][28] ), .G_ik(\g[0][28] ), 
        .P_k1j(\p[0][27] ), .G_k1j(\g[0][27] ), .P_ij(\p[1][13] ), .G_ij_BAR(
        \g[1][13] ) );
  PG_BLOCK_851 Block_Stage_TWO_1 ( .P_ik(\p[1][3] ), .G_ik(\g[1][3] ), .P_k1j(
        1'b0), .G_k1j(\g[1][2] ), .G_ij_BAR(\g[2][1] ) );
  PG_BLOCK_850 Block_Stage_TWO_2 ( .P_ik(\p[1][5] ), .G_ik(\g[1][5] ), .P_k1j(
        \p[1][4] ), .G_k1j(\g[1][4] ), .P_ij(\p[2][2] ), .G_ij(\g[2][2] ) );
  PG_BLOCK_849 Block_Stage_TWO_3 ( .P_ik(\p[1][7] ), .G_ik(\g[1][7] ), .P_k1j(
        \p[1][6] ), .G_k1j(\g[1][6] ), .P_ij(\p[2][3] ), .G_ij(\g[2][3] ) );
  PG_BLOCK_848 Block_Stage_TWO_4 ( .P_ik(\p[1][9] ), .G_ik(\g[1][9] ), .P_k1j(
        \p[1][8] ), .G_k1j(\g[1][8] ), .P_ij(\p[2][4] ), .G_ij(\g[2][4] ) );
  PG_BLOCK_847 Block_Stage_TWO_5 ( .P_ik(\p[1][11] ), .G_ik(\g[1][11] ), 
        .P_k1j(\p[1][10] ), .G_k1j(\g[1][10] ), .P_ij(\p[2][5] ), .G_ij(
        \g[2][5] ) );
  PG_BLOCK_846 Block_Stage_TWO_6 ( .P_ik(\p[1][13] ), .P_k1j(\p[1][12] ), 
        .G_k1j(\g[1][12] ), .P_ij(\p[2][6] ), .G_ij(\g[2][6] ), .G_ik_BAR(
        \g[1][13] ) );
  G_BLOCK_236 g_3 ( .P_ik(1'b0), .G_k1j(1'b0), .G_ij(Cout[2]), .G_ik_BAR(
        \g[2][1] ) );
  PG_BLOCK_836 Block_Stage_THREE_1 ( .P_ik(\p[2][3] ), .G_ik(\g[2][3] ), 
        .P_k1j(\p[2][2] ), .G_k1j(\g[2][2] ), .P_ij(\p[3][1] ), .G_ij(
        \g[3][1] ) );
  PG_BLOCK_835 Block_Stage_THREE_2 ( .P_ik(\p[2][5] ), .G_ik(\g[2][5] ), 
        .P_k1j(\p[2][4] ), .G_k1j(\g[2][4] ), .P_ij(\p[3][2] ), .G_ij(
        \g[3][2] ) );
  G_BLOCK_235 g_4_c12_c16_0 ( .P_ik(\p[2][2] ), .G_ik(\g[2][2] ), .G_k1j(
        Cout[2]), .G_ij(Cout[3]) );
  G_BLOCK_234 g_4_c12_c16_1 ( .P_ik(\p[3][1] ), .G_ik(\g[3][1] ), .G_k1j(
        Cout[2]), .G_ij(Cout[4]) );
  PG_BLOCK_829 Block_stage_FOUR_2_0 ( .P_ik(\p[2][6] ), .G_ik(\g[2][6] ), 
        .P_k1j(\p[3][2] ), .G_k1j(\g[3][2] ), .P_ij(\p[4][2] ), .G_ij(
        \g[4][2] ) );
  G_BLOCK_233 Block_stage_FIVE_4 ( .P_ik(\p[2][4] ), .G_ik(\g[2][4] ), .G_k1j(
        Cout[4]), .G_ij(Cout[5]) );
  G_BLOCK_232 Block_stage_FIVE_5 ( .P_ik(\p[3][2] ), .G_ik(\g[3][2] ), .G_k1j(
        Cout[4]), .G_ij(Cout[6]) );
  G_BLOCK_231 Block_stage_FIVE_6 ( .P_ik(\p[4][2] ), .G_ik(\g[4][2] ), .G_k1j(
        Cout[4]), .G_ij(Cout[7]) );
endmodule


module FA_1792 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1791 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1790 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1789 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_448 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_1792 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_1791 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_1790 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_1789 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_224 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_224 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_448 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0)
         );
  MUX_2to1_N4_224 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_1784 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1783 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1782 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1781 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_446 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1784 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1783 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1782 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1781 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_223 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_223 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_446 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  MUX_2to1_N4_223 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_1776 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1775 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1774 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1773 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_444 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1776 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1775 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1774 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1773 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1772 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_1771 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1770 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1769 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_443 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1772 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1771 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1770 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1769 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_222 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
  MUX2_X1 U2 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U3 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U4 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
endmodule


module carry_select_block_N4_222 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_444 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_443 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_222 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_1768 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1767 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4;

  XOR2_X1 U1 ( .A(Ci), .B(A), .Z(n1) );
  XOR2_X1 U2 ( .A(B), .B(n1), .Z(S) );
  NAND2_X1 U3 ( .A1(B), .A2(Ci), .ZN(n2) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n3) );
  NAND2_X1 U5 ( .A1(Ci), .A2(A), .ZN(n4) );
  NAND3_X1 U6 ( .A1(n2), .A2(n3), .A3(n4), .ZN(Co) );
endmodule


module FA_1766 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1765 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_442 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1768 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1767 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1766 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1765 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1764 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(S) );
endmodule


module FA_1763 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1762 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4, n5;

  XNOR2_X1 U1 ( .A(Ci), .B(n5), .ZN(S) );
  AND2_X1 U2 ( .A1(n1), .A2(n2), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n5) );
  INV_X1 U4 ( .A(B), .ZN(n1) );
  INV_X1 U5 ( .A(A), .ZN(n2) );
  INV_X1 U6 ( .A(Ci), .ZN(n3) );
  OAI22_X1 U7 ( .A1(n3), .A2(n4), .B1(n2), .B2(n1), .ZN(Co) );
endmodule


module FA_1761 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_441 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1764 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1763 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1762 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1761 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_221 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;
  wire   n1, n2, n3;

  NAND2_X1 U1 ( .A1(n1), .A2(n3), .ZN(Y[3]) );
  NAND2_X1 U2 ( .A1(IN0[3]), .A2(n2), .ZN(n1) );
  INV_X1 U3 ( .A(SEL), .ZN(n2) );
  NAND2_X1 U4 ( .A1(IN1[3]), .A2(SEL), .ZN(n3) );
  MUX2_X1 U5 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U6 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U7 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
endmodule


module carry_select_block_N4_221 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_442 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_441 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_221 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_1760 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1759 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1758 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1757 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_440 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1760 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1759 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1758 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1757 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1756 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_1755 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1754 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1753 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_439 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1756 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1755 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1754 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1753 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_220 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X2 U1 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
  MUX2_X1 U2 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U3 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U4 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
endmodule


module carry_select_block_N4_220 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_440 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_439 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_220 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_1752 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1751 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1750 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1749 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_438 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1752 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1751 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1750 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1749 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1748 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_1747 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1746 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1745 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_437 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1748 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1747 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1746 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1745 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_219 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;
  wire   n1, n2, n3;

  NAND2_X1 U1 ( .A1(n3), .A2(n1), .ZN(Y[3]) );
  NAND2_X1 U2 ( .A1(n2), .A2(IN0[3]), .ZN(n1) );
  INV_X1 U3 ( .A(SEL), .ZN(n2) );
  NAND2_X1 U4 ( .A1(IN1[3]), .A2(SEL), .ZN(n3) );
  MUX2_X1 U5 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U6 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U7 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
endmodule


module carry_select_block_N4_219 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_438 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_437 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_219 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_1744 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1743 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1742 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n1) );
  XOR2_X1 U2 ( .A(Ci), .B(n1), .Z(S) );
  NAND2_X1 U3 ( .A1(Ci), .A2(B), .ZN(n2) );
  NAND2_X1 U4 ( .A1(Ci), .A2(A), .ZN(n3) );
  NAND2_X1 U5 ( .A1(B), .A2(A), .ZN(n4) );
  NAND3_X1 U6 ( .A1(n2), .A2(n3), .A3(n4), .ZN(Co) );
endmodule


module FA_1741 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(Ci), .B(n1), .ZN(S) );
endmodule


module RCA_N4_436 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1744 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1743 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1742 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1741 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1740 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_1739 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1738 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(n1) );
  NOR2_X1 U2 ( .A1(B), .A2(A), .ZN(n3) );
  OAI21_X1 U3 ( .B1(n2), .B2(n3), .A(n1), .ZN(Co) );
  INV_X1 U4 ( .A(Ci), .ZN(n2) );
  XOR2_X1 U5 ( .A(B), .B(A), .Z(n4) );
  XOR2_X1 U6 ( .A(Ci), .B(n4), .Z(S) );
endmodule


module FA_1737 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(Ci), .B(n1), .ZN(S) );
endmodule


module RCA_N4_435 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1740 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1739 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1738 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1737 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_218 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X2 U1 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
  MUX2_X1 U2 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U3 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U4 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
endmodule


module carry_select_block_N4_218 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_436 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_435 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_218 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_1736 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(S) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(Co) );
endmodule


module FA_1735 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1734 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1733 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_434 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1736 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1735 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1734 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1733 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1732 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(S) );
  OR2_X1 U2 ( .A1(A), .A2(B), .ZN(Co) );
endmodule


module FA_1731 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1730 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1729 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_433 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1732 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1731 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1730 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1729 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_217 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U2 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U3 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U4 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
endmodule


module carry_select_block_N4_217 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_434 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_433 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_217 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module SUMGENERATOR_Nblocks16_bits_per_block4_14 ( A, B, CARRY_SELECT, SUM );
  input [63:0] A;
  input [63:0] B;
  input [15:0] CARRY_SELECT;
  output [63:0] SUM;


  carry_select_block_N4_224 block_n_1 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(
        B[3:0]), .S(SUM[3:0]), .Ci(1'b0) );
  carry_select_block_N4_223 block_n_2 ( .A(A[7:4]), .B(B[7:4]), .S(SUM[7:4]), 
        .Ci(1'b0) );
  carry_select_block_N4_222 block_n_3 ( .A(A[11:8]), .B(B[11:8]), .S(SUM[11:8]), .Ci(CARRY_SELECT[2]) );
  carry_select_block_N4_221 block_n_4 ( .A(A[15:12]), .B(B[15:12]), .S(
        SUM[15:12]), .Ci(CARRY_SELECT[3]) );
  carry_select_block_N4_220 block_n_5 ( .A(A[19:16]), .B(B[19:16]), .S(
        SUM[19:16]), .Ci(CARRY_SELECT[4]) );
  carry_select_block_N4_219 block_n_6 ( .A(A[23:20]), .B(B[23:20]), .S(
        SUM[23:20]), .Ci(CARRY_SELECT[5]) );
  carry_select_block_N4_218 block_n_7 ( .A(A[27:24]), .B(B[27:24]), .S(
        SUM[27:24]), .Ci(CARRY_SELECT[6]) );
  carry_select_block_N4_217 block_n_8 ( .A(A[31:28]), .B(B[31:28]), .S(
        SUM[31:28]), .Ci(CARRY_SELECT[7]) );
endmodule


module ADDER_P4_N_BIT64_14 ( A, B, add_sub, Cout, SUM );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input add_sub;
  output Cout;
  wire   n1, n2, n4, n5, n6;
  wire   [63:0] B_xor;
  wire   [15:0] tmp_co;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42;
  assign B_xor[31] = B[31];
  assign B_xor[30] = B[30];
  assign B_xor[29] = B[29];
  assign B_xor[28] = B[28];
  assign B_xor[27] = B[27];
  assign B_xor[26] = B[26];
  assign B_xor[25] = B[25];
  assign B_xor[23] = B[23];
  assign B_xor[22] = B[22];
  assign B_xor[21] = B[21];
  assign B_xor[20] = B[20];
  assign B_xor[19] = B[19];
  assign B_xor[18] = B[18];
  assign B_xor[17] = B[17];
  assign B_xor[16] = B[16];
  assign B_xor[15] = B[15];
  assign B_xor[14] = B[14];
  assign B_xor[13] = B[13];
  assign B_xor[12] = B[12];
  assign B_xor[11] = B[11];
  assign B_xor[10] = B[10];
  assign B_xor[9] = B[9];
  assign B_xor[8] = B[8];
  assign B_xor[7] = B[7];
  assign B_xor[6] = B[6];
  assign B_xor[5] = B[5];
  assign B_xor[4] = B[4];
  assign B_xor[3] = B[3];
  assign B_xor[2] = B[2];
  assign B_xor[1] = B[1];
  assign B_xor[0] = B[0];

  CARRY_GENERATOR_Nbit64_14 CLA_SPARSE_TREE ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, A[27:4], 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, B_xor[27:25], B[24], B_xor[23:4], 1'b0, 1'b0, 1'b0, 1'b0}), 
        .Cin(1'b0), .Cout({SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, tmp_co[7:2], SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10}) );
  SUMGENERATOR_Nblocks16_bits_per_block4_14 CSA ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, A[31:4], 1'b0, 1'b0, 1'b0, 1'b0}), .B({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B_xor[31:25], B[24], 
        B_xor[23:16], n1, n6, n2, B_xor[12:8], n4, B_xor[6:0]}), 
        .CARRY_SELECT({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        tmp_co[7:2], 1'b0, 1'b0}), .SUM({SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SUM[31:0]}) );
  BUF_X1 U1 ( .A(B_xor[13]), .Z(n2) );
  BUF_X1 U2 ( .A(B_xor[15]), .Z(n1) );
  CLKBUF_X1 U3 ( .A(B_xor[7]), .Z(n4) );
  INV_X1 U4 ( .A(B_xor[14]), .ZN(n5) );
  INV_X1 U5 ( .A(n5), .ZN(n6) );
endmodule


module PG_NETWORK_826 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_825 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_824 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_823 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_822 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_821 ( op1, op2, g, p );
  input op1, op2;
  output g, p;
  wire   n1;

  XNOR2_X1 U1 ( .A(op2), .B(n1), .ZN(p) );
  INV_X1 U2 ( .A(op1), .ZN(n1) );
  AND2_X1 U3 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_820 ( op1, op2, g, p );
  input op1, op2;
  output g, p;
  wire   n1;

  XNOR2_X1 U1 ( .A(op2), .B(n1), .ZN(p) );
  INV_X1 U2 ( .A(op1), .ZN(n1) );
  AND2_X1 U3 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_819 ( op1, op2, g, p );
  input op1, op2;
  output g, p;
  wire   n1;

  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XNOR2_X1 U2 ( .A(op2), .B(n1), .ZN(p) );
  INV_X1 U3 ( .A(op1), .ZN(n1) );
endmodule


module PG_NETWORK_818 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_817 ( op1, op2, g, p );
  input op1, op2;
  output g, p;
  wire   n1;

  XNOR2_X1 U1 ( .A(op2), .B(n1), .ZN(p) );
  INV_X1 U2 ( .A(op1), .ZN(n1) );
  AND2_X1 U3 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_816 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_815 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_814 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_813 ( op1, op2, g, p );
  input op1, op2;
  output g, p;
  wire   n1;

  XNOR2_X1 U1 ( .A(op2), .B(n1), .ZN(p) );
  INV_X1 U2 ( .A(op1), .ZN(n1) );
  AND2_X1 U3 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_812 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_811 ( op1, op2, g, p );
  input op1, op2;
  output g, p;
  wire   n1;

  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XNOR2_X1 U2 ( .A(op2), .B(n1), .ZN(p) );
  INV_X1 U3 ( .A(op1), .ZN(n1) );
endmodule


module PG_NETWORK_810 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_809 ( op1, op2, g, p );
  input op1, op2;
  output g, p;
  wire   n1;

  XNOR2_X1 U1 ( .A(op2), .B(n1), .ZN(p) );
  INV_X1 U2 ( .A(op1), .ZN(n1) );
  AND2_X1 U3 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_808 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_807 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_806 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_805 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  XOR2_X1 U1 ( .A(op1), .B(op2), .Z(p) );
  AND2_X1 U2 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_BLOCK_817 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij_BAR );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij_BAR;


  AOI21_X1 U1 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(G_ij_BAR) );
endmodule


module PG_BLOCK_816 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_815 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(G_ij) );
  AND2_X1 U2 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U3 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
endmodule


module PG_BLOCK_814 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AOI21_X1 U1 ( .B1(P_ik), .B2(G_k1j), .A(G_ik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(G_ij) );
  AND2_X1 U3 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
endmodule


module PG_BLOCK_813 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1, n2;

  AND2_X1 U1 ( .A1(P_k1j), .A2(P_ik), .ZN(P_ij) );
  NAND2_X1 U2 ( .A1(n2), .A2(n1), .ZN(G_ij) );
  INV_X1 U3 ( .A(G_ik), .ZN(n1) );
  NAND2_X1 U4 ( .A1(P_ik), .A2(G_k1j), .ZN(n2) );
endmodule


module PG_BLOCK_812 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_811 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_810 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AOI21_X1 U1 ( .B1(P_ik), .B2(G_k1j), .A(G_ik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(G_ij) );
  AND2_X1 U3 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
endmodule


module PG_BLOCK_809 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1, n2;

  NAND2_X1 U1 ( .A1(n2), .A2(n1), .ZN(G_ij) );
  INV_X1 U2 ( .A(G_ik), .ZN(n1) );
  NAND2_X1 U3 ( .A1(P_ik), .A2(G_k1j), .ZN(n2) );
  AND2_X1 U4 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
endmodule


module PG_BLOCK_808 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_807 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij_BAR );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij_BAR;


  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(G_k1j), .A(G_ik), .ZN(G_ij_BAR) );
endmodule


module PG_BLOCK_788 ( P_ik, P_k1j, G_k1j, P_ij, G_ij_BAR, G_ik_BAR );
  input P_ik, P_k1j, G_k1j, G_ik_BAR;
  output P_ij, G_ij_BAR;
  wire   G_ik;
  assign G_ij_BAR = G_ik;
  assign G_ik = G_ik_BAR;

endmodule


module PG_BLOCK_787 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AOI21_X1 U1 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(G_ij) );
  AND2_X1 U3 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
endmodule


module PG_BLOCK_786 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1, n2;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  NAND2_X1 U2 ( .A1(G_k1j), .A2(P_ik), .ZN(n1) );
  INV_X1 U3 ( .A(G_ik), .ZN(n2) );
  NAND2_X1 U4 ( .A1(n2), .A2(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_785 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_784 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1, n2;

  NAND2_X1 U1 ( .A1(n2), .A2(n1), .ZN(G_ij) );
  NAND2_X1 U2 ( .A1(G_k1j), .A2(P_ik), .ZN(n1) );
  INV_X1 U3 ( .A(G_ik), .ZN(n2) );
  AND2_X1 U4 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
endmodule


module PG_BLOCK_783 ( P_ik, P_k1j, G_k1j, P_ij, G_ij, G_ik_BAR );
  input P_ik, P_k1j, G_k1j, G_ik_BAR;
  output P_ij, G_ij;
  wire   G_ik, n1;
  assign G_ik = G_ik_BAR;

  NAND2_X1 U1 ( .A1(n1), .A2(G_ik), .ZN(G_ij) );
  NAND2_X1 U2 ( .A1(P_ik), .A2(G_k1j), .ZN(n1) );
  AND2_X1 U3 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
endmodule


module G_BLOCK_219 ( P_ik, G_k1j, G_ij, G_ik_BAR );
  input P_ik, G_k1j, G_ik_BAR;
  output G_ij;
  wire   G_ik;
  assign G_ik = G_ik_BAR;

  INV_X1 U1 ( .A(G_ik), .ZN(G_ij) );
endmodule


module PG_BLOCK_773 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1, n2;

  NAND2_X1 U1 ( .A1(n2), .A2(n1), .ZN(G_ij) );
  NAND2_X1 U2 ( .A1(P_ik), .A2(G_k1j), .ZN(n1) );
  INV_X1 U3 ( .A(G_ik), .ZN(n2) );
  AND2_X1 U4 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
endmodule


module PG_BLOCK_772 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1, n2;

  NAND2_X1 U1 ( .A1(n2), .A2(n1), .ZN(G_ij) );
  NAND2_X1 U2 ( .A1(P_ik), .A2(G_k1j), .ZN(n1) );
  INV_X1 U3 ( .A(G_ik), .ZN(n2) );
  AND2_X1 U4 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
endmodule


module G_BLOCK_218 ( P_ik, G_ik, G_k1j, G_ij );
  input P_ik, G_ik, G_k1j;
  output G_ij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(G_ij) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(G_k1j), .A(G_ik), .ZN(n1) );
endmodule


module G_BLOCK_217 ( P_ik, G_ik, G_k1j, G_ij );
  input P_ik, G_ik, G_k1j;
  output G_ij;
  wire   n1;

  OR2_X2 U1 ( .A1(G_ik), .A2(n1), .ZN(G_ij) );
  AND2_X1 U2 ( .A1(P_ik), .A2(G_k1j), .ZN(n1) );
endmodule


module PG_BLOCK_766 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1, n2;

  NAND2_X1 U1 ( .A1(n2), .A2(n1), .ZN(G_ij) );
  INV_X1 U2 ( .A(G_ik), .ZN(n1) );
  NAND2_X1 U3 ( .A1(G_k1j), .A2(P_ik), .ZN(n2) );
  AND2_X1 U4 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
endmodule


module G_BLOCK_216 ( P_ik, G_ik, G_k1j, G_ij );
  input P_ik, G_ik, G_k1j;
  output G_ij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(G_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
endmodule


module G_BLOCK_215 ( P_ik, G_ik, G_k1j, G_ij );
  input P_ik, G_ik, G_k1j;
  output G_ij;
  wire   n1;

  OR2_X2 U1 ( .A1(n1), .A2(G_ik), .ZN(G_ij) );
  AND2_X1 U2 ( .A1(G_k1j), .A2(P_ik), .ZN(n1) );
endmodule


module G_BLOCK_214 ( P_ik, G_ik, G_k1j, G_ij );
  input P_ik, G_ik, G_k1j;
  output G_ij;
  wire   n2;

  OR2_X1 U1 ( .A1(G_ik), .A2(n2), .ZN(G_ij) );
  AND2_X1 U2 ( .A1(G_k1j), .A2(P_ik), .ZN(n2) );
endmodule


module CARRY_GENERATOR_Nbit64_13 ( A, B, Cin, Cout );
  input [63:0] A;
  input [63:0] B;
  output [16:0] Cout;
  input Cin;
  wire   \p[4][2] , \p[3][2] , \p[3][1] , \p[2][6] , \p[2][5] , \p[2][4] ,
         \p[2][3] , \p[2][2] , \p[1][13] , \p[1][12] , \p[1][11] , \p[1][10] ,
         \p[1][9] , \p[1][8] , \p[1][7] , \p[1][6] , \p[1][5] , \p[1][4] ,
         \p[0][28] , \p[0][27] , \p[0][26] , \p[0][25] , \p[0][24] ,
         \p[0][23] , \p[0][22] , \p[0][21] , \p[0][20] , \p[0][19] ,
         \p[0][18] , \p[0][17] , \p[0][16] , \p[0][15] , \p[0][14] ,
         \p[0][13] , \p[0][12] , \p[0][11] , \p[0][10] , \p[0][9] , \p[0][8] ,
         \g[4][2] , \g[3][2] , \g[3][1] , \g[2][6] , \g[2][5] , \g[2][4] ,
         \g[2][3] , \g[2][2] , \g[2][1] , \g[1][13] , \g[1][12] , \g[1][11] ,
         \g[1][10] , \g[1][9] , \g[1][8] , \g[1][7] , \g[1][6] , \g[1][5] ,
         \g[1][4] , \g[1][3] , \g[0][28] , \g[0][27] , \g[0][26] , \g[0][25] ,
         \g[0][24] , \g[0][23] , \g[0][22] , \g[0][21] , \g[0][20] ,
         \g[0][19] , \g[0][18] , \g[0][17] , \g[0][16] , \g[0][15] ,
         \g[0][14] , \g[0][13] , \g[0][12] , \g[0][11] , \g[0][10] , \g[0][9] ,
         \g[0][8] , \g[0][7] , n1;

  PG_NETWORK_826 Block_PG_NET_7 ( .op1(A[6]), .op2(B[6]), .g(\g[0][7] ) );
  PG_NETWORK_825 Block_PG_NET_8 ( .op1(A[7]), .op2(B[7]), .g(\g[0][8] ), .p(
        \p[0][8] ) );
  PG_NETWORK_824 Block_PG_NET_9 ( .op1(A[8]), .op2(B[8]), .g(\g[0][9] ), .p(
        \p[0][9] ) );
  PG_NETWORK_823 Block_PG_NET_10 ( .op1(A[9]), .op2(B[9]), .g(\g[0][10] ), .p(
        \p[0][10] ) );
  PG_NETWORK_822 Block_PG_NET_11 ( .op1(A[10]), .op2(B[10]), .g(\g[0][11] ), 
        .p(\p[0][11] ) );
  PG_NETWORK_821 Block_PG_NET_12 ( .op1(A[11]), .op2(B[11]), .g(\g[0][12] ), 
        .p(\p[0][12] ) );
  PG_NETWORK_820 Block_PG_NET_13 ( .op1(A[12]), .op2(B[12]), .g(\g[0][13] ), 
        .p(\p[0][13] ) );
  PG_NETWORK_819 Block_PG_NET_14 ( .op1(A[13]), .op2(B[13]), .g(\g[0][14] ), 
        .p(\p[0][14] ) );
  PG_NETWORK_818 Block_PG_NET_15 ( .op1(A[14]), .op2(B[14]), .g(\g[0][15] ), 
        .p(\p[0][15] ) );
  PG_NETWORK_817 Block_PG_NET_16 ( .op1(A[15]), .op2(B[15]), .g(\g[0][16] ), 
        .p(\p[0][16] ) );
  PG_NETWORK_816 Block_PG_NET_17 ( .op1(A[16]), .op2(B[16]), .g(\g[0][17] ), 
        .p(\p[0][17] ) );
  PG_NETWORK_815 Block_PG_NET_18 ( .op1(A[17]), .op2(B[17]), .g(\g[0][18] ), 
        .p(\p[0][18] ) );
  PG_NETWORK_814 Block_PG_NET_19 ( .op1(A[18]), .op2(B[18]), .g(\g[0][19] ), 
        .p(\p[0][19] ) );
  PG_NETWORK_813 Block_PG_NET_20 ( .op1(A[19]), .op2(B[19]), .g(\g[0][20] ), 
        .p(\p[0][20] ) );
  PG_NETWORK_812 Block_PG_NET_21 ( .op1(A[20]), .op2(B[20]), .g(\g[0][21] ), 
        .p(\p[0][21] ) );
  PG_NETWORK_811 Block_PG_NET_22 ( .op1(A[21]), .op2(B[21]), .g(\g[0][22] ), 
        .p(\p[0][22] ) );
  PG_NETWORK_810 Block_PG_NET_23 ( .op1(A[22]), .op2(B[22]), .g(\g[0][23] ), 
        .p(\p[0][23] ) );
  PG_NETWORK_809 Block_PG_NET_24 ( .op1(A[23]), .op2(B[23]), .g(\g[0][24] ), 
        .p(\p[0][24] ) );
  PG_NETWORK_808 Block_PG_NET_25 ( .op1(A[24]), .op2(B[24]), .g(\g[0][25] ), 
        .p(\p[0][25] ) );
  PG_NETWORK_807 Block_PG_NET_26 ( .op1(A[25]), .op2(B[25]), .g(\g[0][26] ), 
        .p(\p[0][26] ) );
  PG_NETWORK_806 Block_PG_NET_27 ( .op1(A[26]), .op2(B[26]), .g(\g[0][27] ), 
        .p(\p[0][27] ) );
  PG_NETWORK_805 Block_PG_NET_28 ( .op1(A[27]), .op2(B[27]), .g(\g[0][28] ), 
        .p(\p[0][28] ) );
  PG_BLOCK_817 Block_Stage_ONE_3 ( .P_ik(\p[0][8] ), .G_ik(\g[0][8] ), .P_k1j(
        1'b0), .G_k1j(\g[0][7] ), .G_ij_BAR(\g[1][3] ) );
  PG_BLOCK_816 Block_Stage_ONE_4 ( .P_ik(\p[0][10] ), .G_ik(\g[0][10] ), 
        .P_k1j(\p[0][9] ), .G_k1j(\g[0][9] ), .P_ij(\p[1][4] ), .G_ij(
        \g[1][4] ) );
  PG_BLOCK_815 Block_Stage_ONE_5 ( .P_ik(\p[0][12] ), .G_ik(\g[0][12] ), 
        .P_k1j(\p[0][11] ), .G_k1j(\g[0][11] ), .P_ij(\p[1][5] ), .G_ij(
        \g[1][5] ) );
  PG_BLOCK_814 Block_Stage_ONE_6 ( .P_ik(\p[0][14] ), .G_ik(\g[0][14] ), 
        .P_k1j(\p[0][13] ), .G_k1j(\g[0][13] ), .P_ij(\p[1][6] ), .G_ij(
        \g[1][6] ) );
  PG_BLOCK_813 Block_Stage_ONE_7 ( .P_ik(\p[0][16] ), .G_ik(\g[0][16] ), 
        .P_k1j(\p[0][15] ), .G_k1j(\g[0][15] ), .P_ij(\p[1][7] ), .G_ij(
        \g[1][7] ) );
  PG_BLOCK_812 Block_Stage_ONE_8 ( .P_ik(\p[0][18] ), .G_ik(\g[0][18] ), 
        .P_k1j(\p[0][17] ), .G_k1j(\g[0][17] ), .P_ij(\p[1][8] ), .G_ij(
        \g[1][8] ) );
  PG_BLOCK_811 Block_Stage_ONE_9 ( .P_ik(\p[0][20] ), .G_ik(\g[0][20] ), 
        .P_k1j(\p[0][19] ), .G_k1j(\g[0][19] ), .P_ij(\p[1][9] ), .G_ij(
        \g[1][9] ) );
  PG_BLOCK_810 Block_Stage_ONE_10 ( .P_ik(\p[0][22] ), .G_ik(\g[0][22] ), 
        .P_k1j(\p[0][21] ), .G_k1j(\g[0][21] ), .P_ij(\p[1][10] ), .G_ij(
        \g[1][10] ) );
  PG_BLOCK_809 Block_Stage_ONE_11 ( .P_ik(\p[0][24] ), .G_ik(\g[0][24] ), 
        .P_k1j(\p[0][23] ), .G_k1j(\g[0][23] ), .P_ij(\p[1][11] ), .G_ij(
        \g[1][11] ) );
  PG_BLOCK_808 Block_Stage_ONE_12 ( .P_ik(\p[0][26] ), .G_ik(\g[0][26] ), 
        .P_k1j(\p[0][25] ), .G_k1j(\g[0][25] ), .P_ij(\p[1][12] ), .G_ij(
        \g[1][12] ) );
  PG_BLOCK_807 Block_Stage_ONE_13 ( .P_ik(\p[0][28] ), .G_ik(\g[0][28] ), 
        .P_k1j(\p[0][27] ), .G_k1j(\g[0][27] ), .P_ij(\p[1][13] ), .G_ij_BAR(
        \g[1][13] ) );
  PG_BLOCK_788 Block_Stage_TWO_1 ( .P_ik(1'b0), .P_k1j(1'b0), .G_k1j(1'b0), 
        .G_ij_BAR(\g[2][1] ), .G_ik_BAR(\g[1][3] ) );
  PG_BLOCK_787 Block_Stage_TWO_2 ( .P_ik(\p[1][5] ), .G_ik(\g[1][5] ), .P_k1j(
        \p[1][4] ), .G_k1j(\g[1][4] ), .P_ij(\p[2][2] ), .G_ij(\g[2][2] ) );
  PG_BLOCK_786 Block_Stage_TWO_3 ( .P_ik(\p[1][7] ), .G_ik(\g[1][7] ), .P_k1j(
        \p[1][6] ), .G_k1j(\g[1][6] ), .P_ij(\p[2][3] ), .G_ij(\g[2][3] ) );
  PG_BLOCK_785 Block_Stage_TWO_4 ( .P_ik(\p[1][9] ), .G_ik(\g[1][9] ), .P_k1j(
        \p[1][8] ), .G_k1j(\g[1][8] ), .P_ij(\p[2][4] ), .G_ij(\g[2][4] ) );
  PG_BLOCK_784 Block_Stage_TWO_5 ( .P_ik(\p[1][11] ), .G_ik(\g[1][11] ), 
        .P_k1j(\p[1][10] ), .G_k1j(\g[1][10] ), .P_ij(\p[2][5] ), .G_ij(
        \g[2][5] ) );
  PG_BLOCK_783 Block_Stage_TWO_6 ( .P_ik(\p[1][13] ), .P_k1j(\p[1][12] ), 
        .G_k1j(\g[1][12] ), .P_ij(\p[2][6] ), .G_ij(\g[2][6] ), .G_ik_BAR(
        \g[1][13] ) );
  G_BLOCK_219 g_3 ( .P_ik(1'b0), .G_k1j(1'b0), .G_ij(Cout[2]), .G_ik_BAR(
        \g[2][1] ) );
  PG_BLOCK_773 Block_Stage_THREE_1 ( .P_ik(\p[2][3] ), .G_ik(\g[2][3] ), 
        .P_k1j(\p[2][2] ), .G_k1j(\g[2][2] ), .P_ij(\p[3][1] ), .G_ij(
        \g[3][1] ) );
  PG_BLOCK_772 Block_Stage_THREE_2 ( .P_ik(\p[2][5] ), .G_ik(\g[2][5] ), 
        .P_k1j(\p[2][4] ), .G_k1j(\g[2][4] ), .P_ij(\p[3][2] ), .G_ij(
        \g[3][2] ) );
  G_BLOCK_218 g_4_c12_c16_0 ( .P_ik(\p[2][2] ), .G_ik(\g[2][2] ), .G_k1j(
        Cout[2]), .G_ij(Cout[3]) );
  G_BLOCK_217 g_4_c12_c16_1 ( .P_ik(\p[3][1] ), .G_ik(\g[3][1] ), .G_k1j(
        Cout[2]), .G_ij(Cout[4]) );
  PG_BLOCK_766 Block_stage_FOUR_2_0 ( .P_ik(\p[2][6] ), .G_ik(\g[2][6] ), 
        .P_k1j(\p[3][2] ), .G_k1j(\g[3][2] ), .P_ij(\p[4][2] ), .G_ij(
        \g[4][2] ) );
  G_BLOCK_216 Block_stage_FIVE_4 ( .P_ik(\p[2][4] ), .G_ik(\g[2][4] ), .G_k1j(
        Cout[4]), .G_ij(Cout[5]) );
  G_BLOCK_215 Block_stage_FIVE_5 ( .P_ik(\p[3][2] ), .G_ik(\g[3][2] ), .G_k1j(
        n1), .G_ij(Cout[6]) );
  G_BLOCK_214 Block_stage_FIVE_6 ( .P_ik(\p[4][2] ), .G_ik(\g[4][2] ), .G_k1j(
        n1), .G_ij(Cout[7]) );
  BUF_X1 U1 ( .A(Cout[4]), .Z(n1) );
endmodule


module FA_1664 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1663 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1662 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1661 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_416 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_1664 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_1663 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_1662 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_1661 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_208 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_208 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_416 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0)
         );
  MUX_2to1_N4_208 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_1656 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1655 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1654 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1653 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_414 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \CTMP[3] ;

  FA_1656 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_1655 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_1654 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(1'b0), .S(S[2]), .Co(\CTMP[3] ) );
  FA_1653 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(\CTMP[3] ), .S(S[3]) );
endmodule


module MUX_2to1_N4_207 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_207 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_414 RCA_0 ( .A({A[3:2], 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0) );
  MUX_2to1_N4_207 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_1648 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1647 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1646 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1645 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_412 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1648 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1647 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1646 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1645 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1644 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_1643 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1642 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1641 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_411 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1644 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1643 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1642 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1641 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_206 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U3 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U4 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
endmodule


module carry_select_block_N4_206 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_412 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_411 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_206 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_1640 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1639 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1638 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1637 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_410 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1640 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1639 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1638 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1637 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1636 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_1635 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1634 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1633 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_409 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1636 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1635 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1634 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1633 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_205 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
  MUX2_X1 U2 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U3 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U4 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
endmodule


module carry_select_block_N4_205 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_410 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_409 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_205 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_1632 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1631 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1630 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1629 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_408 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1632 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1631 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1630 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1629 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1628 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_1627 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1626 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1625 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_407 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1628 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1627 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1626 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1625 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_204 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U3 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U4 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
endmodule


module carry_select_block_N4_204 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_408 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_407 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_204 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_1624 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  BUF_X1 U1 ( .A(B), .Z(n1) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U3 ( .A(n1), .B(A), .Z(S) );
endmodule


module FA_1623 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1622 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1621 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(Ci), .B(n1), .ZN(S) );
endmodule


module RCA_N4_406 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1624 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1623 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1622 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1621 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1620 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  BUF_X1 U1 ( .A(B), .Z(n1) );
  OR2_X1 U2 ( .A1(B), .A2(A), .ZN(Co) );
  XNOR2_X1 U3 ( .A(n1), .B(A), .ZN(S) );
endmodule


module FA_1619 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1618 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4;

  OAI21_X1 U1 ( .B1(n2), .B2(n1), .A(n4), .ZN(Co) );
  NOR2_X1 U2 ( .A1(B), .A2(A), .ZN(n1) );
  INV_X1 U3 ( .A(Ci), .ZN(n2) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n3) );
  XOR2_X1 U5 ( .A(Ci), .B(n3), .Z(S) );
  NAND2_X1 U6 ( .A1(B), .A2(A), .ZN(n4) );
endmodule


module FA_1617 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(Ci), .B(n1), .ZN(S) );
endmodule


module RCA_N4_405 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1620 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1619 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1618 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1617 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_203 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X2 U1 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
  MUX2_X1 U2 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U3 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U4 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
endmodule


module carry_select_block_N4_203 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_406 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_405 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_203 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_1616 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1615 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1614 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1613 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_404 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1616 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1615 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1614 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1613 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1612 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(S) );
endmodule


module FA_1611 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1610 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1609 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(Ci), .B(n1), .ZN(S) );
endmodule


module RCA_N4_403 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1612 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1611 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1610 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1609 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_202 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
  MUX2_X1 U3 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U4 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
endmodule


module carry_select_block_N4_202 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_404 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_403 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_202 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_1608 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1607 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1606 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1605 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_402 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1608 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1607 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1606 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1605 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1604 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(S) );
endmodule


module FA_1603 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1602 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1601 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_401 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1604 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1603 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1602 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1601 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_201 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;
  wire   n1;

  MUX2_X1 U1 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U2 ( .A(IN0[2]), .B(IN1[2]), .S(n1), .Z(Y[2]) );
  MUX2_X1 U3 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  BUF_X1 U4 ( .A(SEL), .Z(n1) );
  MUX2_X1 U5 ( .A(IN0[3]), .B(IN1[3]), .S(n1), .Z(Y[3]) );
endmodule


module carry_select_block_N4_201 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_402 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_401 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_201 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module SUMGENERATOR_Nblocks16_bits_per_block4_13 ( A, B, CARRY_SELECT, SUM );
  input [63:0] A;
  input [63:0] B;
  input [15:0] CARRY_SELECT;
  output [63:0] SUM;


  carry_select_block_N4_208 block_n_1 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(
        B[3:0]), .S(SUM[3:0]), .Ci(1'b0) );
  carry_select_block_N4_207 block_n_2 ( .A({A[7:6], 1'b0, 1'b0}), .B(B[7:4]), 
        .S(SUM[7:4]), .Ci(1'b0) );
  carry_select_block_N4_206 block_n_3 ( .A(A[11:8]), .B(B[11:8]), .S(SUM[11:8]), .Ci(CARRY_SELECT[2]) );
  carry_select_block_N4_205 block_n_4 ( .A(A[15:12]), .B(B[15:12]), .S(
        SUM[15:12]), .Ci(CARRY_SELECT[3]) );
  carry_select_block_N4_204 block_n_5 ( .A(A[19:16]), .B(B[19:16]), .S(
        SUM[19:16]), .Ci(CARRY_SELECT[4]) );
  carry_select_block_N4_203 block_n_6 ( .A(A[23:20]), .B(B[23:20]), .S(
        SUM[23:20]), .Ci(CARRY_SELECT[5]) );
  carry_select_block_N4_202 block_n_7 ( .A(A[27:24]), .B(B[27:24]), .S(
        SUM[27:24]), .Ci(CARRY_SELECT[6]) );
  carry_select_block_N4_201 block_n_8 ( .A(A[31:28]), .B(B[31:28]), .S(
        SUM[31:28]), .Ci(CARRY_SELECT[7]) );
endmodule


module ADDER_P4_N_BIT64_13 ( A, B, add_sub, Cout, SUM );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input add_sub;
  output Cout;
  wire   n1, n2, n3, n4;
  wire   [63:0] B_xor;
  wire   [15:0] tmp_co;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42;
  assign B_xor[31] = B[31];
  assign B_xor[30] = B[30];
  assign B_xor[29] = B[29];
  assign B_xor[28] = B[28];
  assign B_xor[27] = B[27];
  assign B_xor[26] = B[26];
  assign B_xor[25] = B[25];
  assign B_xor[24] = B[24];
  assign B_xor[23] = B[23];
  assign B_xor[22] = B[22];
  assign B_xor[21] = B[21];
  assign B_xor[20] = B[20];
  assign B_xor[19] = B[19];
  assign B_xor[18] = B[18];
  assign B_xor[17] = B[17];
  assign B_xor[16] = B[16];
  assign B_xor[15] = B[15];
  assign B_xor[14] = B[14];
  assign B_xor[13] = B[13];
  assign B_xor[12] = B[12];
  assign B_xor[11] = B[11];
  assign B_xor[10] = B[10];
  assign B_xor[9] = B[9];
  assign B_xor[8] = B[8];
  assign B_xor[7] = B[7];
  assign B_xor[6] = B[6];
  assign B_xor[5] = B[5];
  assign B_xor[4] = B[4];
  assign B_xor[3] = B[3];
  assign B_xor[2] = B[2];
  assign B_xor[1] = B[1];
  assign B_xor[0] = B[0];

  CARRY_GENERATOR_Nbit64_13 CLA_SPARSE_TREE ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, A[27:6], 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, B_xor[27:6], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .Cin(1'b0), .Cout({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, tmp_co[7:2], 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10}) );
  SUMGENERATOR_Nblocks16_bits_per_block4_13 CSA ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, A[31:6], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B_xor[31:24], n2, 
        B_xor[22:16], n4, B_xor[14], n1, B_xor[12], n3, B_xor[10:0]}), 
        .CARRY_SELECT({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        tmp_co[7:2], 1'b0, 1'b0}), .SUM({SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SUM[31:0]}) );
  BUF_X1 U1 ( .A(B_xor[13]), .Z(n1) );
  BUF_X1 U2 ( .A(B_xor[23]), .Z(n2) );
  BUF_X1 U3 ( .A(B_xor[11]), .Z(n3) );
  BUF_X1 U4 ( .A(B_xor[15]), .Z(n4) );
endmodule


module PG_NETWORK_760 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_759 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_758 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_757 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_756 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_755 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_754 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_753 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_752 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_751 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_750 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_749 ( op1, op2, g, p );
  input op1, op2;
  output g, p;
  wire   n1;

  XNOR2_X1 U1 ( .A(op2), .B(n1), .ZN(p) );
  INV_X1 U2 ( .A(op1), .ZN(n1) );
  AND2_X1 U3 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_748 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_747 ( op1, op2, g, p );
  input op1, op2;
  output g, p;
  wire   n1;

  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XNOR2_X1 U2 ( .A(op2), .B(n1), .ZN(p) );
  INV_X1 U3 ( .A(op1), .ZN(n1) );
endmodule


module PG_NETWORK_746 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_745 ( op1, op2, g, p );
  input op1, op2;
  output g, p;
  wire   n1;

  XNOR2_X1 U1 ( .A(op2), .B(n1), .ZN(p) );
  INV_X1 U2 ( .A(op1), .ZN(n1) );
  AND2_X1 U3 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_744 ( op1, op2, g, p );
  input op1, op2;
  output g, p;
  wire   n1;

  XNOR2_X1 U1 ( .A(op2), .B(n1), .ZN(p) );
  INV_X1 U2 ( .A(op1), .ZN(n1) );
  AND2_X1 U3 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_743 ( op1, op2, g, p );
  input op1, op2;
  output g, p;
  wire   n1;

  XNOR2_X1 U1 ( .A(op2), .B(n1), .ZN(p) );
  INV_X1 U2 ( .A(op1), .ZN(n1) );
  AND2_X1 U3 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_742 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  XOR2_X1 U1 ( .A(op1), .B(op2), .Z(p) );
  AND2_X1 U2 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_741 ( op1, op2, g, p );
  input op1, op2;
  output g, p;
  wire   n1;

  XNOR2_X1 U1 ( .A(op2), .B(n1), .ZN(p) );
  INV_X1 U2 ( .A(op1), .ZN(n1) );
  AND2_X1 U3 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_BLOCK_753 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AOI21_X1 U1 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_752 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_751 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_750 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(G_k1j), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_749 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_748 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(G_k1j), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_747 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AOI21_X1 U1 ( .B1(P_ik), .B2(G_k1j), .A(G_ik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(G_ij) );
  AND2_X1 U3 ( .A1(P_k1j), .A2(P_ik), .ZN(P_ij) );
endmodule


module PG_BLOCK_746 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1, n2;

  NAND2_X1 U1 ( .A1(n2), .A2(n1), .ZN(G_ij) );
  INV_X1 U2 ( .A(G_ik), .ZN(n1) );
  NAND2_X1 U3 ( .A1(P_ik), .A2(G_k1j), .ZN(n2) );
  AND2_X1 U4 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
endmodule


module PG_BLOCK_745 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1, n2;

  NAND2_X1 U1 ( .A1(n2), .A2(n1), .ZN(G_ij) );
  INV_X1 U2 ( .A(G_ik), .ZN(n1) );
  NAND2_X1 U3 ( .A1(P_ik), .A2(G_k1j), .ZN(n2) );
  AND2_X1 U4 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
endmodule


module PG_BLOCK_744 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1, n2;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  NAND2_X1 U2 ( .A1(n2), .A2(n1), .ZN(G_ij) );
  INV_X1 U3 ( .A(G_ik), .ZN(n1) );
  NAND2_X1 U4 ( .A1(P_ik), .A2(G_k1j), .ZN(n2) );
endmodule


module PG_BLOCK_724 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij_BAR );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij_BAR;


  AOI21_X1 U1 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(G_ij_BAR) );
endmodule


module PG_BLOCK_723 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_722 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n2;

  OR2_X1 U1 ( .A1(n2), .A2(G_ik), .ZN(G_ij) );
  AND2_X1 U2 ( .A1(G_k1j), .A2(P_ik), .ZN(n2) );
  AND2_X1 U3 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
endmodule


module PG_BLOCK_721 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1, n2;

  NAND2_X1 U1 ( .A1(n1), .A2(n2), .ZN(G_ij) );
  INV_X1 U2 ( .A(G_ik), .ZN(n1) );
  NAND2_X1 U3 ( .A1(G_k1j), .A2(P_ik), .ZN(n2) );
  AND2_X1 U4 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
endmodule


module PG_BLOCK_720 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1, n2;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  NAND2_X1 U2 ( .A1(n1), .A2(n2), .ZN(G_ij) );
  INV_X1 U3 ( .A(G_ik), .ZN(n1) );
  NAND2_X1 U4 ( .A1(P_ik), .A2(G_k1j), .ZN(n2) );
endmodule


module PG_BLOCK_710 ( P_ik, G_ik, P_k1j, P_ij, G_ij_BAR, G_k1j_BAR );
  input P_ik, G_ik, P_k1j, G_k1j_BAR;
  output P_ij, G_ij_BAR;
  wire   G_k1j, n1, n3;
  assign G_k1j = G_k1j_BAR;

  NOR2_X1 U1 ( .A1(G_ik), .A2(n1), .ZN(G_ij_BAR) );
  AND2_X1 U2 ( .A1(P_ik), .A2(n3), .ZN(n1) );
  INV_X1 U3 ( .A(G_k1j), .ZN(n3) );
endmodule


module PG_BLOCK_709 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1, n2;

  NAND2_X1 U1 ( .A1(n2), .A2(n1), .ZN(G_ij) );
  NAND2_X1 U2 ( .A1(P_ik), .A2(G_k1j), .ZN(n1) );
  INV_X1 U3 ( .A(G_ik), .ZN(n2) );
  AND2_X1 U4 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
endmodule


module G_BLOCK_201 ( P_ik, G_k1j, G_ij, G_ik_BAR );
  input P_ik, G_k1j, G_ik_BAR;
  output G_ij;
  wire   G_ik;
  assign G_ik = G_ik_BAR;

  INV_X1 U1 ( .A(G_ik), .ZN(G_ij) );
endmodule


module G_BLOCK_200 ( P_ik, G_k1j, G_ij, G_ik_BAR );
  input P_ik, G_k1j, G_ik_BAR;
  output G_ij;
  wire   G_ik;
  assign G_ik = G_ik_BAR;

  INV_X1 U1 ( .A(G_ik), .ZN(G_ij) );
endmodule


module PG_BLOCK_703 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1, n2;

  NAND2_X1 U1 ( .A1(n1), .A2(n2), .ZN(G_ij) );
  NAND2_X1 U2 ( .A1(G_k1j), .A2(P_ik), .ZN(n1) );
  INV_X1 U3 ( .A(G_ik), .ZN(n2) );
  AND2_X1 U4 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
endmodule


module G_BLOCK_199 ( P_ik, G_ik, G_k1j, G_ij );
  input P_ik, G_ik, G_k1j;
  output G_ij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(G_ij) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(G_k1j), .A(G_ik), .ZN(n1) );
endmodule


module G_BLOCK_198 ( P_ik, G_ik, G_k1j, G_ij );
  input P_ik, G_ik, G_k1j;
  output G_ij;
  wire   n1;

  AOI21_X1 U1 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(G_ij) );
endmodule


module G_BLOCK_197 ( P_ik, G_ik, G_k1j, G_ij );
  input P_ik, G_ik, G_k1j;
  output G_ij;
  wire   n1;

  OR2_X2 U1 ( .A1(G_ik), .A2(n1), .ZN(G_ij) );
  AND2_X1 U2 ( .A1(P_ik), .A2(G_k1j), .ZN(n1) );
endmodule


module CARRY_GENERATOR_Nbit64_12 ( A, B, Cin, Cout );
  input [63:0] A;
  input [63:0] B;
  output [16:0] Cout;
  input Cin;
  wire   \p[4][2] , \p[3][2] , \p[2][6] , \p[2][5] , \p[2][4] , \p[2][3] ,
         \p[1][13] , \p[1][12] , \p[1][11] , \p[1][10] , \p[1][9] , \p[1][8] ,
         \p[1][7] , \p[1][6] , \p[1][5] , \p[0][28] , \p[0][27] , \p[0][26] ,
         \p[0][25] , \p[0][24] , \p[0][23] , \p[0][22] , \p[0][21] ,
         \p[0][20] , \p[0][19] , \p[0][18] , \p[0][17] , \p[0][16] ,
         \p[0][15] , \p[0][14] , \p[0][13] , \p[0][12] , \p[0][11] ,
         \p[0][10] , \g[4][2] , \g[3][2] , \g[3][1] , \g[2][6] , \g[2][5] ,
         \g[2][4] , \g[2][3] , \g[2][2] , \g[1][13] , \g[1][12] , \g[1][11] ,
         \g[1][10] , \g[1][9] , \g[1][8] , \g[1][7] , \g[1][6] , \g[1][5] ,
         \g[1][4] , \g[0][28] , \g[0][27] , \g[0][26] , \g[0][25] , \g[0][24] ,
         \g[0][23] , \g[0][22] , \g[0][21] , \g[0][20] , \g[0][19] ,
         \g[0][18] , \g[0][17] , \g[0][16] , \g[0][15] , \g[0][14] ,
         \g[0][13] , \g[0][12] , \g[0][11] , \g[0][10] , \g[0][9] ;

  PG_NETWORK_760 Block_PG_NET_9 ( .op1(A[8]), .op2(B[8]), .g(\g[0][9] ) );
  PG_NETWORK_759 Block_PG_NET_10 ( .op1(A[9]), .op2(B[9]), .g(\g[0][10] ), .p(
        \p[0][10] ) );
  PG_NETWORK_758 Block_PG_NET_11 ( .op1(A[10]), .op2(B[10]), .g(\g[0][11] ), 
        .p(\p[0][11] ) );
  PG_NETWORK_757 Block_PG_NET_12 ( .op1(A[11]), .op2(B[11]), .g(\g[0][12] ), 
        .p(\p[0][12] ) );
  PG_NETWORK_756 Block_PG_NET_13 ( .op1(A[12]), .op2(B[12]), .g(\g[0][13] ), 
        .p(\p[0][13] ) );
  PG_NETWORK_755 Block_PG_NET_14 ( .op1(A[13]), .op2(B[13]), .g(\g[0][14] ), 
        .p(\p[0][14] ) );
  PG_NETWORK_754 Block_PG_NET_15 ( .op1(A[14]), .op2(B[14]), .g(\g[0][15] ), 
        .p(\p[0][15] ) );
  PG_NETWORK_753 Block_PG_NET_16 ( .op1(A[15]), .op2(B[15]), .g(\g[0][16] ), 
        .p(\p[0][16] ) );
  PG_NETWORK_752 Block_PG_NET_17 ( .op1(A[16]), .op2(B[16]), .g(\g[0][17] ), 
        .p(\p[0][17] ) );
  PG_NETWORK_751 Block_PG_NET_18 ( .op1(A[17]), .op2(B[17]), .g(\g[0][18] ), 
        .p(\p[0][18] ) );
  PG_NETWORK_750 Block_PG_NET_19 ( .op1(A[18]), .op2(B[18]), .g(\g[0][19] ), 
        .p(\p[0][19] ) );
  PG_NETWORK_749 Block_PG_NET_20 ( .op1(A[19]), .op2(B[19]), .g(\g[0][20] ), 
        .p(\p[0][20] ) );
  PG_NETWORK_748 Block_PG_NET_21 ( .op1(A[20]), .op2(B[20]), .g(\g[0][21] ), 
        .p(\p[0][21] ) );
  PG_NETWORK_747 Block_PG_NET_22 ( .op1(A[21]), .op2(B[21]), .g(\g[0][22] ), 
        .p(\p[0][22] ) );
  PG_NETWORK_746 Block_PG_NET_23 ( .op1(A[22]), .op2(B[22]), .g(\g[0][23] ), 
        .p(\p[0][23] ) );
  PG_NETWORK_745 Block_PG_NET_24 ( .op1(A[23]), .op2(B[23]), .g(\g[0][24] ), 
        .p(\p[0][24] ) );
  PG_NETWORK_744 Block_PG_NET_25 ( .op1(A[24]), .op2(B[24]), .g(\g[0][25] ), 
        .p(\p[0][25] ) );
  PG_NETWORK_743 Block_PG_NET_26 ( .op1(A[25]), .op2(B[25]), .g(\g[0][26] ), 
        .p(\p[0][26] ) );
  PG_NETWORK_742 Block_PG_NET_27 ( .op1(A[26]), .op2(B[26]), .g(\g[0][27] ), 
        .p(\p[0][27] ) );
  PG_NETWORK_741 Block_PG_NET_28 ( .op1(A[27]), .op2(B[27]), .g(\g[0][28] ), 
        .p(\p[0][28] ) );
  PG_BLOCK_753 Block_Stage_ONE_4 ( .P_ik(\p[0][10] ), .G_ik(\g[0][10] ), 
        .P_k1j(1'b0), .G_k1j(\g[0][9] ), .G_ij(\g[1][4] ) );
  PG_BLOCK_752 Block_Stage_ONE_5 ( .P_ik(\p[0][12] ), .G_ik(\g[0][12] ), 
        .P_k1j(\p[0][11] ), .G_k1j(\g[0][11] ), .P_ij(\p[1][5] ), .G_ij(
        \g[1][5] ) );
  PG_BLOCK_751 Block_Stage_ONE_6 ( .P_ik(\p[0][14] ), .G_ik(\g[0][14] ), 
        .P_k1j(\p[0][13] ), .G_k1j(\g[0][13] ), .P_ij(\p[1][6] ), .G_ij(
        \g[1][6] ) );
  PG_BLOCK_750 Block_Stage_ONE_7 ( .P_ik(\p[0][16] ), .G_ik(\g[0][16] ), 
        .P_k1j(\p[0][15] ), .G_k1j(\g[0][15] ), .P_ij(\p[1][7] ), .G_ij(
        \g[1][7] ) );
  PG_BLOCK_749 Block_Stage_ONE_8 ( .P_ik(\p[0][18] ), .G_ik(\g[0][18] ), 
        .P_k1j(\p[0][17] ), .G_k1j(\g[0][17] ), .P_ij(\p[1][8] ), .G_ij(
        \g[1][8] ) );
  PG_BLOCK_748 Block_Stage_ONE_9 ( .P_ik(\p[0][20] ), .G_ik(\g[0][20] ), 
        .P_k1j(\p[0][19] ), .G_k1j(\g[0][19] ), .P_ij(\p[1][9] ), .G_ij(
        \g[1][9] ) );
  PG_BLOCK_747 Block_Stage_ONE_10 ( .P_ik(\p[0][22] ), .G_ik(\g[0][22] ), 
        .P_k1j(\p[0][21] ), .G_k1j(\g[0][21] ), .P_ij(\p[1][10] ), .G_ij(
        \g[1][10] ) );
  PG_BLOCK_746 Block_Stage_ONE_11 ( .P_ik(\p[0][24] ), .G_ik(\g[0][24] ), 
        .P_k1j(\p[0][23] ), .G_k1j(\g[0][23] ), .P_ij(\p[1][11] ), .G_ij(
        \g[1][11] ) );
  PG_BLOCK_745 Block_Stage_ONE_12 ( .P_ik(\p[0][26] ), .G_ik(\g[0][26] ), 
        .P_k1j(\p[0][25] ), .G_k1j(\g[0][25] ), .P_ij(\p[1][12] ), .G_ij(
        \g[1][12] ) );
  PG_BLOCK_744 Block_Stage_ONE_13 ( .P_ik(\p[0][28] ), .G_ik(\g[0][28] ), 
        .P_k1j(\p[0][27] ), .G_k1j(\g[0][27] ), .P_ij(\p[1][13] ), .G_ij(
        \g[1][13] ) );
  PG_BLOCK_724 Block_Stage_TWO_2 ( .P_ik(\p[1][5] ), .G_ik(\g[1][5] ), .P_k1j(
        1'b0), .G_k1j(\g[1][4] ), .G_ij_BAR(\g[2][2] ) );
  PG_BLOCK_723 Block_Stage_TWO_3 ( .P_ik(\p[1][7] ), .G_ik(\g[1][7] ), .P_k1j(
        \p[1][6] ), .G_k1j(\g[1][6] ), .P_ij(\p[2][3] ), .G_ij(\g[2][3] ) );
  PG_BLOCK_722 Block_Stage_TWO_4 ( .P_ik(\p[1][9] ), .G_ik(\g[1][9] ), .P_k1j(
        \p[1][8] ), .G_k1j(\g[1][8] ), .P_ij(\p[2][4] ), .G_ij(\g[2][4] ) );
  PG_BLOCK_721 Block_Stage_TWO_5 ( .P_ik(\p[1][11] ), .G_ik(\g[1][11] ), 
        .P_k1j(\p[1][10] ), .G_k1j(\g[1][10] ), .P_ij(\p[2][5] ), .G_ij(
        \g[2][5] ) );
  PG_BLOCK_720 Block_Stage_TWO_6 ( .P_ik(\p[1][13] ), .G_ik(\g[1][13] ), 
        .P_k1j(\p[1][12] ), .G_k1j(\g[1][12] ), .P_ij(\p[2][6] ), .G_ij(
        \g[2][6] ) );
  PG_BLOCK_710 Block_Stage_THREE_1 ( .P_ik(\p[2][3] ), .G_ik(\g[2][3] ), 
        .P_k1j(1'b0), .G_ij_BAR(\g[3][1] ), .G_k1j_BAR(\g[2][2] ) );
  PG_BLOCK_709 Block_Stage_THREE_2 ( .P_ik(\p[2][5] ), .G_ik(\g[2][5] ), 
        .P_k1j(\p[2][4] ), .G_k1j(\g[2][4] ), .P_ij(\p[3][2] ), .G_ij(
        \g[3][2] ) );
  G_BLOCK_201 g_4_c12_c16_0 ( .P_ik(1'b0), .G_k1j(1'b0), .G_ij(Cout[3]), 
        .G_ik_BAR(\g[2][2] ) );
  G_BLOCK_200 g_4_c12_c16_1 ( .P_ik(1'b0), .G_k1j(1'b0), .G_ij(Cout[4]), 
        .G_ik_BAR(\g[3][1] ) );
  PG_BLOCK_703 Block_stage_FOUR_2_0 ( .P_ik(\p[2][6] ), .G_ik(\g[2][6] ), 
        .P_k1j(\p[3][2] ), .G_k1j(\g[3][2] ), .P_ij(\p[4][2] ), .G_ij(
        \g[4][2] ) );
  G_BLOCK_199 Block_stage_FIVE_4 ( .P_ik(\p[2][4] ), .G_ik(\g[2][4] ), .G_k1j(
        Cout[4]), .G_ij(Cout[5]) );
  G_BLOCK_198 Block_stage_FIVE_5 ( .P_ik(\p[3][2] ), .G_ik(\g[3][2] ), .G_k1j(
        Cout[4]), .G_ij(Cout[6]) );
  G_BLOCK_197 Block_stage_FIVE_6 ( .P_ik(\p[4][2] ), .G_ik(\g[4][2] ), .G_k1j(
        Cout[4]), .G_ij(Cout[7]) );
endmodule


module FA_1536 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1535 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1534 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1533 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_384 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_1536 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_1535 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_1534 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_1533 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_192 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_192 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_384 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0)
         );
  MUX_2to1_N4_192 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_1528 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1527 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1526 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1525 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_382 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_1528 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_1527 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_1526 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_1525 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_191 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_191 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_382 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0)
         );
  MUX_2to1_N4_191 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_1520 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1519 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1518 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1517 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_380 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1520 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1519 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1518 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1517 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_190 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_190 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_380 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  MUX_2to1_N4_190 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_1512 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1511 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1510 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1509 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n2) );
  XNOR2_X1 U2 ( .A(n2), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_378 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1512 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1511 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1510 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1509 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1508 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_1507 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1506 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1505 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n2) );
  XNOR2_X1 U2 ( .A(n2), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_377 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1508 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1507 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1506 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1505 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_189 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U3 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U4 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
endmodule


module carry_select_block_N4_189 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_378 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_377 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_189 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_1504 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1503 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1502 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1501 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_376 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1504 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1503 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1502 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1501 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1500 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_1499 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1498 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1497 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_375 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1500 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1499 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1498 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1497 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_188 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U3 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U4 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
endmodule


module carry_select_block_N4_188 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_376 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_375 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_188 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_1496 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1495 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1494 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1493 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_374 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1496 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1495 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1494 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1493 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1492 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_1491 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1490 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1489 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_373 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1492 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1491 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1490 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1489 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_187 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U3 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U4 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
endmodule


module carry_select_block_N4_187 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_374 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_373 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_187 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_1488 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1487 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1486 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1485 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_372 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1488 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1487 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1486 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1485 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1484 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  BUF_X1 U1 ( .A(B), .Z(n1) );
  OR2_X1 U2 ( .A1(B), .A2(A), .ZN(Co) );
  XNOR2_X1 U3 ( .A(A), .B(n1), .ZN(S) );
endmodule


module FA_1483 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1482 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1481 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(Ci), .B(n1), .ZN(S) );
endmodule


module RCA_N4_371 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1484 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1483 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1482 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1481 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_186 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;
  wire   n1, n2, n3;

  NAND2_X1 U1 ( .A1(n3), .A2(n1), .ZN(Y[3]) );
  NAND2_X1 U2 ( .A1(IN0[3]), .A2(n2), .ZN(n1) );
  INV_X1 U3 ( .A(SEL), .ZN(n2) );
  NAND2_X1 U4 ( .A1(IN1[3]), .A2(SEL), .ZN(n3) );
  MUX2_X1 U5 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U6 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U7 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
endmodule


module carry_select_block_N4_186 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_372 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_371 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_186 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_1480 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1479 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4;

  OAI21_X1 U1 ( .B1(B), .B2(Ci), .A(A), .ZN(n1) );
  OAI21_X1 U2 ( .B1(n2), .B2(n3), .A(n1), .ZN(Co) );
  INV_X1 U3 ( .A(B), .ZN(n2) );
  INV_X1 U4 ( .A(Ci), .ZN(n3) );
  XOR2_X1 U5 ( .A(B), .B(A), .Z(n4) );
  XOR2_X1 U6 ( .A(Ci), .B(n4), .Z(S) );
endmodule


module FA_1478 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4;

  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(n2) );
  OR2_X1 U2 ( .A1(B), .A2(A), .ZN(n3) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n4) );
  NAND2_X1 U4 ( .A1(n1), .A2(n2), .ZN(Co) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n3), .ZN(n1) );
  XNOR2_X1 U6 ( .A(Ci), .B(n4), .ZN(S) );
endmodule


module FA_1477 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(Ci), .B(n1), .ZN(S) );
endmodule


module RCA_N4_370 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1480 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1479 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1478 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1477 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1476 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(S) );
endmodule


module FA_1475 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4;

  NAND2_X1 U1 ( .A1(n1), .A2(n4), .ZN(Co) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n2), .ZN(n1) );
  OR2_X1 U3 ( .A1(B), .A2(A), .ZN(n2) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n3) );
  XOR2_X1 U5 ( .A(Ci), .B(n3), .Z(S) );
  NAND2_X1 U6 ( .A1(B), .A2(A), .ZN(n4) );
endmodule


module FA_1474 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4;

  OR2_X1 U1 ( .A1(B), .A2(A), .ZN(n3) );
  NAND2_X1 U2 ( .A1(B), .A2(A), .ZN(n1) );
  NAND2_X1 U3 ( .A1(n2), .A2(n1), .ZN(Co) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n2) );
  XOR2_X1 U5 ( .A(B), .B(A), .Z(n4) );
  XOR2_X1 U6 ( .A(Ci), .B(n4), .Z(S) );
endmodule


module FA_1473 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(Ci), .B(n1), .ZN(S) );
endmodule


module RCA_N4_369 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1476 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1475 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1474 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1473 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_185 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U3 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U4 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
endmodule


module carry_select_block_N4_185 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_370 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_369 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_185 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module SUMGENERATOR_Nblocks16_bits_per_block4_12 ( A, B, CARRY_SELECT, SUM );
  input [63:0] A;
  input [63:0] B;
  input [15:0] CARRY_SELECT;
  output [63:0] SUM;


  carry_select_block_N4_192 block_n_1 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(
        B[3:0]), .S(SUM[3:0]), .Ci(1'b0) );
  carry_select_block_N4_191 block_n_2 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(
        B[7:4]), .S(SUM[7:4]), .Ci(1'b0) );
  carry_select_block_N4_190 block_n_3 ( .A(A[11:8]), .B(B[11:8]), .S(SUM[11:8]), .Ci(1'b0) );
  carry_select_block_N4_189 block_n_4 ( .A(A[15:12]), .B(B[15:12]), .S(
        SUM[15:12]), .Ci(CARRY_SELECT[3]) );
  carry_select_block_N4_188 block_n_5 ( .A(A[19:16]), .B(B[19:16]), .S(
        SUM[19:16]), .Ci(CARRY_SELECT[4]) );
  carry_select_block_N4_187 block_n_6 ( .A(A[23:20]), .B(B[23:20]), .S(
        SUM[23:20]), .Ci(CARRY_SELECT[5]) );
  carry_select_block_N4_186 block_n_7 ( .A(A[27:24]), .B(B[27:24]), .S(
        SUM[27:24]), .Ci(CARRY_SELECT[6]) );
  carry_select_block_N4_185 block_n_8 ( .A(A[31:28]), .B(B[31:28]), .S(
        SUM[31:28]), .Ci(CARRY_SELECT[7]) );
endmodule


module ADDER_P4_N_BIT64_12 ( A, B, add_sub, Cout, SUM );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input add_sub;
  output Cout;
  wire   n1, n2, n3, n4, n5, n7, n8, n9, n10;
  wire   [63:0] B_xor;
  wire   [15:0] tmp_co;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43;
  assign B_xor[31] = B[31];
  assign B_xor[30] = B[30];
  assign B_xor[29] = B[29];
  assign B_xor[28] = B[28];
  assign B_xor[27] = B[27];
  assign B_xor[26] = B[26];
  assign B_xor[25] = B[25];
  assign B_xor[24] = B[24];
  assign B_xor[23] = B[23];
  assign B_xor[22] = B[22];
  assign B_xor[21] = B[21];
  assign B_xor[20] = B[20];
  assign B_xor[19] = B[19];
  assign B_xor[18] = B[18];
  assign B_xor[17] = B[17];
  assign B_xor[16] = B[16];
  assign B_xor[14] = B[14];
  assign B_xor[13] = B[13];
  assign B_xor[12] = B[12];
  assign B_xor[11] = B[11];
  assign B_xor[10] = B[10];
  assign B_xor[9] = B[9];
  assign B_xor[8] = B[8];
  assign B_xor[7] = B[7];
  assign B_xor[6] = B[6];
  assign B_xor[5] = B[5];
  assign B_xor[4] = B[4];
  assign B_xor[3] = B[3];
  assign B_xor[2] = B[2];
  assign B_xor[1] = B[1];
  assign B_xor[0] = B[0];

  CARRY_GENERATOR_Nbit64_12 CLA_SPARSE_TREE ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, A[27:8], 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B_xor[27:16], B[15], B_xor[14:8], 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Cin(1'b0), .Cout({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, tmp_co[7:3], SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11}) );
  SUMGENERATOR_Nblocks16_bits_per_block4_12 CSA ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, A[31:8], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        B_xor[31:28], n5, n2, n3, B_xor[24], n10, n8, n9, n1, B_xor[19:16], 
        B[15], B_xor[14:0]}), .CARRY_SELECT({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, tmp_co[7:3], 1'b0, 1'b0, 1'b0}), .SUM({
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, SUM[31:0]}) );
  BUF_X1 U1 ( .A(B_xor[25]), .Z(n3) );
  BUF_X1 U2 ( .A(B_xor[26]), .Z(n2) );
  BUF_X1 U3 ( .A(B_xor[20]), .Z(n1) );
  INV_X1 U4 ( .A(B_xor[27]), .ZN(n4) );
  INV_X1 U5 ( .A(n4), .ZN(n5) );
  CLKBUF_X1 U6 ( .A(B_xor[21]), .Z(n9) );
  INV_X1 U7 ( .A(B_xor[22]), .ZN(n7) );
  INV_X1 U8 ( .A(n7), .ZN(n8) );
  BUF_X1 U9 ( .A(B_xor[23]), .Z(n10) );
endmodule


module PG_NETWORK_694 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_693 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_692 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_691 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op1), .A2(op2), .ZN(g) );
  XOR2_X1 U2 ( .A(op1), .B(op2), .Z(p) );
endmodule


module PG_NETWORK_690 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_689 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op1), .A2(op2), .ZN(g) );
  XOR2_X1 U2 ( .A(op1), .B(op2), .Z(p) );
endmodule


module PG_NETWORK_688 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_687 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_686 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_685 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_684 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_683 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_682 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_681 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  XOR2_X1 U1 ( .A(op2), .B(op1), .Z(p) );
  AND2_X1 U2 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_680 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_679 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_678 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_677 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_BLOCK_689 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij_BAR );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij_BAR;


  AOI21_X1 U1 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(G_ij_BAR) );
endmodule


module PG_BLOCK_688 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_687 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(G_k1j), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_686 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_685 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_684 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_683 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij_BAR );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij_BAR;


  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(G_k1j), .A(G_ik), .ZN(G_ij_BAR) );
endmodule


module PG_BLOCK_682 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_681 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_661 ( P_ik, P_k1j, G_k1j, P_ij, G_ij_BAR, G_ik_BAR );
  input P_ik, P_k1j, G_k1j, G_ik_BAR;
  output P_ij, G_ij_BAR;
  wire   G_ik;
  assign G_ij_BAR = G_ik;
  assign G_ik = G_ik_BAR;

endmodule


module PG_BLOCK_660 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_659 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_658 ( P_ik, P_k1j, G_k1j, P_ij, G_ij, G_ik_BAR );
  input P_ik, P_k1j, G_k1j, G_ik_BAR;
  output P_ij, G_ij;
  wire   G_ik, n1;
  assign G_ik = G_ik_BAR;

  NAND2_X1 U1 ( .A1(n1), .A2(G_ik), .ZN(G_ij) );
  NAND2_X1 U2 ( .A1(G_k1j), .A2(P_ik), .ZN(n1) );
  AND2_X1 U3 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
endmodule


module PG_BLOCK_657 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_647 ( P_ik, G_ik, P_k1j, P_ij, G_ij_BAR, G_k1j_BAR );
  input P_ik, G_ik, P_k1j, G_k1j_BAR;
  output P_ij, G_ij_BAR;
  wire   G_k1j, n1;
  assign G_k1j = G_k1j_BAR;

  INV_X1 U1 ( .A(G_k1j), .ZN(n1) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(n1), .A(G_ik), .ZN(G_ij_BAR) );
endmodule


module PG_BLOCK_646 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module G_BLOCK_184 ( P_ik, G_k1j, G_ij, G_ik_BAR );
  input P_ik, G_k1j, G_ik_BAR;
  output G_ij;
  wire   G_ik;
  assign G_ik = G_ik_BAR;

  INV_X1 U1 ( .A(G_ik), .ZN(G_ij) );
endmodule


module G_BLOCK_183 ( P_ik, G_k1j, G_ij, G_ik_BAR );
  input P_ik, G_k1j, G_ik_BAR;
  output G_ij;
  wire   G_ik;
  assign G_ik = G_ik_BAR;

  INV_X1 U1 ( .A(G_ik), .ZN(G_ij) );
endmodule


module PG_BLOCK_640 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module G_BLOCK_182 ( P_ik, G_ik, G_k1j, G_ij );
  input P_ik, G_ik, G_k1j;
  output G_ij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(G_ij) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(G_k1j), .A(G_ik), .ZN(n1) );
endmodule


module G_BLOCK_181 ( P_ik, G_ik, G_k1j, G_ij );
  input P_ik, G_ik, G_k1j;
  output G_ij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(G_ij) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(G_k1j), .A(G_ik), .ZN(n1) );
endmodule


module G_BLOCK_180 ( P_ik, G_ik, G_k1j, G_ij );
  input P_ik, G_ik, G_k1j;
  output G_ij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(G_ij) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(G_k1j), .A(G_ik), .ZN(n1) );
endmodule


module CARRY_GENERATOR_Nbit64_11 ( A, B, Cin, Cout );
  input [63:0] A;
  input [63:0] B;
  output [16:0] Cout;
  input Cin;
  wire   \p[4][2] , \p[3][2] , \p[2][6] , \p[2][5] , \p[2][4] , \p[2][3] ,
         \p[1][13] , \p[1][12] , \p[1][11] , \p[1][10] , \p[1][9] , \p[1][8] ,
         \p[1][7] , \p[1][6] , \p[0][28] , \p[0][27] , \p[0][26] , \p[0][25] ,
         \p[0][24] , \p[0][23] , \p[0][22] , \p[0][21] , \p[0][20] ,
         \p[0][19] , \p[0][18] , \p[0][17] , \p[0][16] , \p[0][15] ,
         \p[0][14] , \p[0][13] , \p[0][12] , \g[4][2] , \g[3][2] , \g[3][1] ,
         \g[2][6] , \g[2][5] , \g[2][4] , \g[2][3] , \g[2][2] , \g[1][13] ,
         \g[1][12] , \g[1][11] , \g[1][10] , \g[1][9] , \g[1][8] , \g[1][7] ,
         \g[1][6] , \g[1][5] , \g[0][28] , \g[0][27] , \g[0][26] , \g[0][25] ,
         \g[0][24] , \g[0][23] , \g[0][22] , \g[0][21] , \g[0][20] ,
         \g[0][19] , \g[0][18] , \g[0][17] , \g[0][16] , \g[0][15] ,
         \g[0][14] , \g[0][13] , \g[0][12] , \g[0][11] ;

  PG_NETWORK_694 Block_PG_NET_11 ( .op1(A[10]), .op2(B[10]), .g(\g[0][11] ) );
  PG_NETWORK_693 Block_PG_NET_12 ( .op1(A[11]), .op2(B[11]), .g(\g[0][12] ), 
        .p(\p[0][12] ) );
  PG_NETWORK_692 Block_PG_NET_13 ( .op1(A[12]), .op2(B[12]), .g(\g[0][13] ), 
        .p(\p[0][13] ) );
  PG_NETWORK_691 Block_PG_NET_14 ( .op1(A[13]), .op2(B[13]), .g(\g[0][14] ), 
        .p(\p[0][14] ) );
  PG_NETWORK_690 Block_PG_NET_15 ( .op1(A[14]), .op2(B[14]), .g(\g[0][15] ), 
        .p(\p[0][15] ) );
  PG_NETWORK_689 Block_PG_NET_16 ( .op1(A[15]), .op2(B[15]), .g(\g[0][16] ), 
        .p(\p[0][16] ) );
  PG_NETWORK_688 Block_PG_NET_17 ( .op1(A[16]), .op2(B[16]), .g(\g[0][17] ), 
        .p(\p[0][17] ) );
  PG_NETWORK_687 Block_PG_NET_18 ( .op1(A[17]), .op2(B[17]), .g(\g[0][18] ), 
        .p(\p[0][18] ) );
  PG_NETWORK_686 Block_PG_NET_19 ( .op1(A[18]), .op2(B[18]), .g(\g[0][19] ), 
        .p(\p[0][19] ) );
  PG_NETWORK_685 Block_PG_NET_20 ( .op1(A[19]), .op2(B[19]), .g(\g[0][20] ), 
        .p(\p[0][20] ) );
  PG_NETWORK_684 Block_PG_NET_21 ( .op1(A[20]), .op2(B[20]), .g(\g[0][21] ), 
        .p(\p[0][21] ) );
  PG_NETWORK_683 Block_PG_NET_22 ( .op1(A[21]), .op2(B[21]), .g(\g[0][22] ), 
        .p(\p[0][22] ) );
  PG_NETWORK_682 Block_PG_NET_23 ( .op1(A[22]), .op2(B[22]), .g(\g[0][23] ), 
        .p(\p[0][23] ) );
  PG_NETWORK_681 Block_PG_NET_24 ( .op1(A[23]), .op2(B[23]), .g(\g[0][24] ), 
        .p(\p[0][24] ) );
  PG_NETWORK_680 Block_PG_NET_25 ( .op1(A[24]), .op2(B[24]), .g(\g[0][25] ), 
        .p(\p[0][25] ) );
  PG_NETWORK_679 Block_PG_NET_26 ( .op1(A[25]), .op2(B[25]), .g(\g[0][26] ), 
        .p(\p[0][26] ) );
  PG_NETWORK_678 Block_PG_NET_27 ( .op1(A[26]), .op2(B[26]), .g(\g[0][27] ), 
        .p(\p[0][27] ) );
  PG_NETWORK_677 Block_PG_NET_28 ( .op1(A[27]), .op2(B[27]), .g(\g[0][28] ), 
        .p(\p[0][28] ) );
  PG_BLOCK_689 Block_Stage_ONE_5 ( .P_ik(\p[0][12] ), .G_ik(\g[0][12] ), 
        .P_k1j(1'b0), .G_k1j(\g[0][11] ), .G_ij_BAR(\g[1][5] ) );
  PG_BLOCK_688 Block_Stage_ONE_6 ( .P_ik(\p[0][14] ), .G_ik(\g[0][14] ), 
        .P_k1j(\p[0][13] ), .G_k1j(\g[0][13] ), .P_ij(\p[1][6] ), .G_ij(
        \g[1][6] ) );
  PG_BLOCK_687 Block_Stage_ONE_7 ( .P_ik(\p[0][16] ), .G_ik(\g[0][16] ), 
        .P_k1j(\p[0][15] ), .G_k1j(\g[0][15] ), .P_ij(\p[1][7] ), .G_ij(
        \g[1][7] ) );
  PG_BLOCK_686 Block_Stage_ONE_8 ( .P_ik(\p[0][18] ), .G_ik(\g[0][18] ), 
        .P_k1j(\p[0][17] ), .G_k1j(\g[0][17] ), .P_ij(\p[1][8] ), .G_ij(
        \g[1][8] ) );
  PG_BLOCK_685 Block_Stage_ONE_9 ( .P_ik(\p[0][20] ), .G_ik(\g[0][20] ), 
        .P_k1j(\p[0][19] ), .G_k1j(\g[0][19] ), .P_ij(\p[1][9] ), .G_ij(
        \g[1][9] ) );
  PG_BLOCK_684 Block_Stage_ONE_10 ( .P_ik(\p[0][22] ), .G_ik(\g[0][22] ), 
        .P_k1j(\p[0][21] ), .G_k1j(\g[0][21] ), .P_ij(\p[1][10] ), .G_ij(
        \g[1][10] ) );
  PG_BLOCK_683 Block_Stage_ONE_11 ( .P_ik(\p[0][24] ), .G_ik(\g[0][24] ), 
        .P_k1j(\p[0][23] ), .G_k1j(\g[0][23] ), .P_ij(\p[1][11] ), .G_ij_BAR(
        \g[1][11] ) );
  PG_BLOCK_682 Block_Stage_ONE_12 ( .P_ik(\p[0][26] ), .G_ik(\g[0][26] ), 
        .P_k1j(\p[0][25] ), .G_k1j(\g[0][25] ), .P_ij(\p[1][12] ), .G_ij(
        \g[1][12] ) );
  PG_BLOCK_681 Block_Stage_ONE_13 ( .P_ik(\p[0][28] ), .G_ik(\g[0][28] ), 
        .P_k1j(\p[0][27] ), .G_k1j(\g[0][27] ), .P_ij(\p[1][13] ), .G_ij(
        \g[1][13] ) );
  PG_BLOCK_661 Block_Stage_TWO_2 ( .P_ik(1'b0), .P_k1j(1'b0), .G_k1j(1'b0), 
        .G_ij_BAR(\g[2][2] ), .G_ik_BAR(\g[1][5] ) );
  PG_BLOCK_660 Block_Stage_TWO_3 ( .P_ik(\p[1][7] ), .G_ik(\g[1][7] ), .P_k1j(
        \p[1][6] ), .G_k1j(\g[1][6] ), .P_ij(\p[2][3] ), .G_ij(\g[2][3] ) );
  PG_BLOCK_659 Block_Stage_TWO_4 ( .P_ik(\p[1][9] ), .G_ik(\g[1][9] ), .P_k1j(
        \p[1][8] ), .G_k1j(\g[1][8] ), .P_ij(\p[2][4] ), .G_ij(\g[2][4] ) );
  PG_BLOCK_658 Block_Stage_TWO_5 ( .P_ik(\p[1][11] ), .P_k1j(\p[1][10] ), 
        .G_k1j(\g[1][10] ), .P_ij(\p[2][5] ), .G_ij(\g[2][5] ), .G_ik_BAR(
        \g[1][11] ) );
  PG_BLOCK_657 Block_Stage_TWO_6 ( .P_ik(\p[1][13] ), .G_ik(\g[1][13] ), 
        .P_k1j(\p[1][12] ), .G_k1j(\g[1][12] ), .P_ij(\p[2][6] ), .G_ij(
        \g[2][6] ) );
  PG_BLOCK_647 Block_Stage_THREE_1 ( .P_ik(\p[2][3] ), .G_ik(\g[2][3] ), 
        .P_k1j(1'b0), .G_ij_BAR(\g[3][1] ), .G_k1j_BAR(\g[2][2] ) );
  PG_BLOCK_646 Block_Stage_THREE_2 ( .P_ik(\p[2][5] ), .G_ik(\g[2][5] ), 
        .P_k1j(\p[2][4] ), .G_k1j(\g[2][4] ), .P_ij(\p[3][2] ), .G_ij(
        \g[3][2] ) );
  G_BLOCK_184 g_4_c12_c16_0 ( .P_ik(1'b0), .G_k1j(1'b0), .G_ij(Cout[3]), 
        .G_ik_BAR(\g[2][2] ) );
  G_BLOCK_183 g_4_c12_c16_1 ( .P_ik(1'b0), .G_k1j(1'b0), .G_ij(Cout[4]), 
        .G_ik_BAR(\g[3][1] ) );
  PG_BLOCK_640 Block_stage_FOUR_2_0 ( .P_ik(\p[2][6] ), .G_ik(\g[2][6] ), 
        .P_k1j(\p[3][2] ), .G_k1j(\g[3][2] ), .P_ij(\p[4][2] ), .G_ij(
        \g[4][2] ) );
  G_BLOCK_182 Block_stage_FIVE_4 ( .P_ik(\p[2][4] ), .G_ik(\g[2][4] ), .G_k1j(
        Cout[4]), .G_ij(Cout[5]) );
  G_BLOCK_181 Block_stage_FIVE_5 ( .P_ik(\p[3][2] ), .G_ik(\g[3][2] ), .G_k1j(
        Cout[4]), .G_ij(Cout[6]) );
  G_BLOCK_180 Block_stage_FIVE_6 ( .P_ik(\p[4][2] ), .G_ik(\g[4][2] ), .G_k1j(
        Cout[4]), .G_ij(Cout[7]) );
endmodule


module FA_1408 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1407 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1406 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1405 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_352 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_1408 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_1407 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_1406 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_1405 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_176 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_176 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_352 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0)
         );
  MUX_2to1_N4_176 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_1400 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1399 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1398 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1397 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_350 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_1400 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_1399 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_1398 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_1397 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_175 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_175 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_350 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0)
         );
  MUX_2to1_N4_175 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_1392 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1391 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1390 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1389 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_348 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \CTMP[3] ;

  FA_1392 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_1391 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_1390 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(1'b0), .S(S[2]), .Co(\CTMP[3] ) );
  FA_1389 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(\CTMP[3] ), .S(S[3]) );
endmodule


module MUX_2to1_N4_174 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_174 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_348 RCA_0 ( .A({A[3:2], 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0) );
  MUX_2to1_N4_174 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_1384 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1383 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1382 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1381 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_346 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1384 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1383 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1382 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1381 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1380 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_1379 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1378 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1377 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_345 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1380 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1379 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1378 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1377 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_173 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U3 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U4 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
endmodule


module carry_select_block_N4_173 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_346 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_345 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_173 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_1376 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1375 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1374 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1373 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_344 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1376 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1375 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1374 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1373 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1372 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_1371 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1370 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1369 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_343 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1372 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1371 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1370 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1369 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_172 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;
  wire   n1;

  BUF_X1 U1 ( .A(SEL), .Z(n1) );
  MUX2_X1 U2 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U3 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U4 ( .A(IN0[2]), .B(IN1[2]), .S(n1), .Z(Y[2]) );
  MUX2_X1 U5 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
endmodule


module carry_select_block_N4_172 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_344 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_343 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_172 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_1368 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1367 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1366 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1365 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_342 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1368 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1367 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1366 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1365 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1364 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_1363 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1362 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1361 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(Ci), .B(n1), .ZN(S) );
endmodule


module RCA_N4_341 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1364 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1363 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1362 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1361 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_171 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U3 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U4 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
endmodule


module carry_select_block_N4_171 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_342 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_341 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_171 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_1360 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1359 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1358 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1357 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_340 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1360 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1359 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1358 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1357 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1356 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_1355 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1354 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1353 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_339 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1356 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1355 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1354 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1353 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_170 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U3 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U4 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
endmodule


module carry_select_block_N4_170 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_340 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_339 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_170 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_1352 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1351 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1350 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1349 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_338 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1352 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1351 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1350 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1349 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1348 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_1347 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1346 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1345 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_337 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1348 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1347 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1346 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1345 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_169 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U3 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U4 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
endmodule


module carry_select_block_N4_169 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_338 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_337 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_169 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module SUMGENERATOR_Nblocks16_bits_per_block4_11 ( A, B, CARRY_SELECT, SUM );
  input [63:0] A;
  input [63:0] B;
  input [15:0] CARRY_SELECT;
  output [63:0] SUM;


  carry_select_block_N4_176 block_n_1 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(
        B[3:0]), .S(SUM[3:0]), .Ci(1'b0) );
  carry_select_block_N4_175 block_n_2 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(
        B[7:4]), .S(SUM[7:4]), .Ci(1'b0) );
  carry_select_block_N4_174 block_n_3 ( .A({A[11:10], 1'b0, 1'b0}), .B(B[11:8]), .S(SUM[11:8]), .Ci(1'b0) );
  carry_select_block_N4_173 block_n_4 ( .A(A[15:12]), .B(B[15:12]), .S(
        SUM[15:12]), .Ci(CARRY_SELECT[3]) );
  carry_select_block_N4_172 block_n_5 ( .A(A[19:16]), .B(B[19:16]), .S(
        SUM[19:16]), .Ci(CARRY_SELECT[4]) );
  carry_select_block_N4_171 block_n_6 ( .A(A[23:20]), .B(B[23:20]), .S(
        SUM[23:20]), .Ci(CARRY_SELECT[5]) );
  carry_select_block_N4_170 block_n_7 ( .A(A[27:24]), .B(B[27:24]), .S(
        SUM[27:24]), .Ci(CARRY_SELECT[6]) );
  carry_select_block_N4_169 block_n_8 ( .A(A[31:28]), .B(B[31:28]), .S(
        SUM[31:28]), .Ci(CARRY_SELECT[7]) );
endmodule


module ADDER_P4_N_BIT64_11 ( A, B, add_sub, Cout, SUM );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input add_sub;
  output Cout;
  wire   n3, n4;
  wire   [63:0] B_xor;
  wire   [15:0] tmp_co;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43;
  assign B_xor[31] = B[31];
  assign B_xor[30] = B[30];
  assign B_xor[29] = B[29];
  assign B_xor[28] = B[28];
  assign B_xor[27] = B[27];
  assign B_xor[26] = B[26];
  assign B_xor[25] = B[25];
  assign B_xor[24] = B[24];
  assign B_xor[23] = B[23];
  assign B_xor[22] = B[22];
  assign B_xor[21] = B[21];
  assign B_xor[20] = B[20];
  assign B_xor[19] = B[19];
  assign B_xor[18] = B[18];
  assign B_xor[17] = B[17];
  assign B_xor[16] = B[16];
  assign B_xor[15] = B[15];
  assign B_xor[14] = B[14];
  assign B_xor[13] = B[13];
  assign B_xor[12] = B[12];
  assign B_xor[11] = B[11];
  assign B_xor[10] = B[10];
  assign B_xor[9] = B[9];
  assign B_xor[8] = B[8];
  assign B_xor[7] = B[7];
  assign B_xor[6] = B[6];
  assign B_xor[5] = B[5];
  assign B_xor[4] = B[4];
  assign B_xor[3] = B[3];
  assign B_xor[2] = B[2];
  assign B_xor[1] = B[1];
  assign B_xor[0] = B[0];

  CARRY_GENERATOR_Nbit64_11 CLA_SPARSE_TREE ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, A[27:10], 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B_xor[27:10], 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Cin(1'b0), 
        .Cout({SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, tmp_co[7:3], SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11}) );
  SUMGENERATOR_Nblocks16_bits_per_block4_11 CSA ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, A[31:16], n4, A[14], n3, A[12:10], 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B_xor[31:0]}), .CARRY_SELECT({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, tmp_co[7:3], 1'b0, 1'b0, 1'b0}), 
        .SUM({SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, SUM[31:0]}) );
  BUF_X1 U1 ( .A(A[13]), .Z(n3) );
  BUF_X1 U2 ( .A(A[15]), .Z(n4) );
endmodule


module PG_NETWORK_628 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_627 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_626 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_625 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  XOR2_X1 U1 ( .A(op1), .B(op2), .Z(p) );
  AND2_X1 U2 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_624 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_623 ( op1, op2, g, p );
  input op1, op2;
  output g, p;
  wire   n1;

  XNOR2_X1 U1 ( .A(op2), .B(n1), .ZN(p) );
  INV_X1 U2 ( .A(op1), .ZN(n1) );
  AND2_X1 U3 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_622 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_621 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_620 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_619 ( op1, op2, g, p );
  input op1, op2;
  output g, p;
  wire   n1;

  XNOR2_X1 U1 ( .A(op2), .B(n1), .ZN(p) );
  INV_X1 U2 ( .A(op1), .ZN(n1) );
  AND2_X1 U3 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_618 ( op1, op2, g, p );
  input op1, op2;
  output g, p;
  wire   n1;

  XNOR2_X1 U1 ( .A(op2), .B(n1), .ZN(p) );
  INV_X1 U2 ( .A(op1), .ZN(n1) );
  AND2_X1 U3 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_617 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_616 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_615 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_614 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_613 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_BLOCK_625 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AOI21_X1 U1 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_624 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_623 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_622 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_621 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(G_k1j), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_620 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij_BAR );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij_BAR;


  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(G_k1j), .A(G_ik), .ZN(G_ij_BAR) );
endmodule


module PG_BLOCK_619 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_618 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_597 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij_BAR );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij_BAR;


  AOI21_X1 U1 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(G_ij_BAR) );
endmodule


module PG_BLOCK_596 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_595 ( P_ik, P_k1j, G_k1j, P_ij, G_ij, G_ik_BAR );
  input P_ik, P_k1j, G_k1j, G_ik_BAR;
  output P_ij, G_ij;
  wire   G_ik, n1;
  assign G_ik = G_ik_BAR;

  NAND2_X1 U1 ( .A1(n1), .A2(G_ik), .ZN(G_ij) );
  NAND2_X1 U2 ( .A1(G_k1j), .A2(P_ik), .ZN(n1) );
  AND2_X1 U3 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
endmodule


module PG_BLOCK_594 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_584 ( P_ik, P_k1j, G_k1j, P_ij, G_ij_BAR, G_ik_BAR );
  input P_ik, P_k1j, G_k1j, G_ik_BAR;
  output P_ij, G_ij_BAR;
  wire   G_ik;
  assign G_ij_BAR = G_ik;
  assign G_ik = G_ik_BAR;

endmodule


module PG_BLOCK_583 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1, n2;

  NAND2_X1 U1 ( .A1(n2), .A2(n1), .ZN(G_ij) );
  NAND2_X1 U2 ( .A1(P_ik), .A2(G_k1j), .ZN(n1) );
  INV_X1 U3 ( .A(G_ik), .ZN(n2) );
  AND2_X1 U4 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
endmodule


module G_BLOCK_166 ( P_ik, G_k1j, G_ij, G_ik_BAR );
  input P_ik, G_k1j, G_ik_BAR;
  output G_ij;
  wire   G_ik;
  assign G_ik = G_ik_BAR;

  INV_X1 U1 ( .A(G_ik), .ZN(G_ij) );
endmodule


module PG_BLOCK_577 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module G_BLOCK_165 ( P_ik, G_ik, G_k1j, G_ij );
  input P_ik, G_ik, G_k1j;
  output G_ij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(G_ij) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(G_k1j), .A(G_ik), .ZN(n1) );
endmodule


module G_BLOCK_164 ( P_ik, G_ik, G_k1j, G_ij );
  input P_ik, G_ik, G_k1j;
  output G_ij;
  wire   n1;

  OR2_X2 U1 ( .A1(G_ik), .A2(n1), .ZN(G_ij) );
  AND2_X1 U2 ( .A1(P_ik), .A2(G_k1j), .ZN(n1) );
endmodule


module G_BLOCK_163 ( P_ik, G_ik, G_k1j, G_ij );
  input P_ik, G_ik, G_k1j;
  output G_ij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(G_ij) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(G_k1j), .A(G_ik), .ZN(n1) );
endmodule


module CARRY_GENERATOR_Nbit64_10 ( A, B, Cin, Cout );
  input [63:0] A;
  input [63:0] B;
  output [16:0] Cout;
  input Cin;
  wire   \p[4][2] , \p[3][2] , \p[2][6] , \p[2][5] , \p[2][4] , \p[1][13] ,
         \p[1][12] , \p[1][11] , \p[1][10] , \p[1][9] , \p[1][8] , \p[1][7] ,
         \p[0][28] , \p[0][27] , \p[0][26] , \p[0][25] , \p[0][24] ,
         \p[0][23] , \p[0][22] , \p[0][21] , \p[0][20] , \p[0][19] ,
         \p[0][18] , \p[0][17] , \p[0][16] , \p[0][15] , \p[0][14] , \g[4][2] ,
         \g[3][2] , \g[3][1] , \g[2][6] , \g[2][5] , \g[2][4] , \g[2][3] ,
         \g[1][13] , \g[1][12] , \g[1][11] , \g[1][10] , \g[1][9] , \g[1][8] ,
         \g[1][7] , \g[1][6] , \g[0][28] , \g[0][27] , \g[0][26] , \g[0][25] ,
         \g[0][24] , \g[0][23] , \g[0][22] , \g[0][21] , \g[0][20] ,
         \g[0][19] , \g[0][18] , \g[0][17] , \g[0][16] , \g[0][15] ,
         \g[0][14] , \g[0][13] ;

  PG_NETWORK_628 Block_PG_NET_13 ( .op1(A[12]), .op2(B[12]), .g(\g[0][13] ) );
  PG_NETWORK_627 Block_PG_NET_14 ( .op1(A[13]), .op2(B[13]), .g(\g[0][14] ), 
        .p(\p[0][14] ) );
  PG_NETWORK_626 Block_PG_NET_15 ( .op1(A[14]), .op2(B[14]), .g(\g[0][15] ), 
        .p(\p[0][15] ) );
  PG_NETWORK_625 Block_PG_NET_16 ( .op1(A[15]), .op2(B[15]), .g(\g[0][16] ), 
        .p(\p[0][16] ) );
  PG_NETWORK_624 Block_PG_NET_17 ( .op1(A[16]), .op2(B[16]), .g(\g[0][17] ), 
        .p(\p[0][17] ) );
  PG_NETWORK_623 Block_PG_NET_18 ( .op1(A[17]), .op2(B[17]), .g(\g[0][18] ), 
        .p(\p[0][18] ) );
  PG_NETWORK_622 Block_PG_NET_19 ( .op1(A[18]), .op2(B[18]), .g(\g[0][19] ), 
        .p(\p[0][19] ) );
  PG_NETWORK_621 Block_PG_NET_20 ( .op1(A[19]), .op2(B[19]), .g(\g[0][20] ), 
        .p(\p[0][20] ) );
  PG_NETWORK_620 Block_PG_NET_21 ( .op1(A[20]), .op2(B[20]), .g(\g[0][21] ), 
        .p(\p[0][21] ) );
  PG_NETWORK_619 Block_PG_NET_22 ( .op1(A[21]), .op2(B[21]), .g(\g[0][22] ), 
        .p(\p[0][22] ) );
  PG_NETWORK_618 Block_PG_NET_23 ( .op1(A[22]), .op2(B[22]), .g(\g[0][23] ), 
        .p(\p[0][23] ) );
  PG_NETWORK_617 Block_PG_NET_24 ( .op1(A[23]), .op2(B[23]), .g(\g[0][24] ), 
        .p(\p[0][24] ) );
  PG_NETWORK_616 Block_PG_NET_25 ( .op1(A[24]), .op2(B[24]), .g(\g[0][25] ), 
        .p(\p[0][25] ) );
  PG_NETWORK_615 Block_PG_NET_26 ( .op1(A[25]), .op2(B[25]), .g(\g[0][26] ), 
        .p(\p[0][26] ) );
  PG_NETWORK_614 Block_PG_NET_27 ( .op1(A[26]), .op2(B[26]), .g(\g[0][27] ), 
        .p(\p[0][27] ) );
  PG_NETWORK_613 Block_PG_NET_28 ( .op1(A[27]), .op2(B[27]), .g(\g[0][28] ), 
        .p(\p[0][28] ) );
  PG_BLOCK_625 Block_Stage_ONE_6 ( .P_ik(\p[0][14] ), .G_ik(\g[0][14] ), 
        .P_k1j(1'b0), .G_k1j(\g[0][13] ), .G_ij(\g[1][6] ) );
  PG_BLOCK_624 Block_Stage_ONE_7 ( .P_ik(\p[0][16] ), .G_ik(\g[0][16] ), 
        .P_k1j(\p[0][15] ), .G_k1j(\g[0][15] ), .P_ij(\p[1][7] ), .G_ij(
        \g[1][7] ) );
  PG_BLOCK_623 Block_Stage_ONE_8 ( .P_ik(\p[0][18] ), .G_ik(\g[0][18] ), 
        .P_k1j(\p[0][17] ), .G_k1j(\g[0][17] ), .P_ij(\p[1][8] ), .G_ij(
        \g[1][8] ) );
  PG_BLOCK_622 Block_Stage_ONE_9 ( .P_ik(\p[0][20] ), .G_ik(\g[0][20] ), 
        .P_k1j(\p[0][19] ), .G_k1j(\g[0][19] ), .P_ij(\p[1][9] ), .G_ij(
        \g[1][9] ) );
  PG_BLOCK_621 Block_Stage_ONE_10 ( .P_ik(\p[0][22] ), .G_ik(\g[0][22] ), 
        .P_k1j(\p[0][21] ), .G_k1j(\g[0][21] ), .P_ij(\p[1][10] ), .G_ij(
        \g[1][10] ) );
  PG_BLOCK_620 Block_Stage_ONE_11 ( .P_ik(\p[0][24] ), .G_ik(\g[0][24] ), 
        .P_k1j(\p[0][23] ), .G_k1j(\g[0][23] ), .P_ij(\p[1][11] ), .G_ij_BAR(
        \g[1][11] ) );
  PG_BLOCK_619 Block_Stage_ONE_12 ( .P_ik(\p[0][26] ), .G_ik(\g[0][26] ), 
        .P_k1j(\p[0][25] ), .G_k1j(\g[0][25] ), .P_ij(\p[1][12] ), .G_ij(
        \g[1][12] ) );
  PG_BLOCK_618 Block_Stage_ONE_13 ( .P_ik(\p[0][28] ), .G_ik(\g[0][28] ), 
        .P_k1j(\p[0][27] ), .G_k1j(\g[0][27] ), .P_ij(\p[1][13] ), .G_ij(
        \g[1][13] ) );
  PG_BLOCK_597 Block_Stage_TWO_3 ( .P_ik(\p[1][7] ), .G_ik(\g[1][7] ), .P_k1j(
        1'b0), .G_k1j(\g[1][6] ), .G_ij_BAR(\g[2][3] ) );
  PG_BLOCK_596 Block_Stage_TWO_4 ( .P_ik(\p[1][9] ), .G_ik(\g[1][9] ), .P_k1j(
        \p[1][8] ), .G_k1j(\g[1][8] ), .P_ij(\p[2][4] ), .G_ij(\g[2][4] ) );
  PG_BLOCK_595 Block_Stage_TWO_5 ( .P_ik(\p[1][11] ), .P_k1j(\p[1][10] ), 
        .G_k1j(\g[1][10] ), .P_ij(\p[2][5] ), .G_ij(\g[2][5] ), .G_ik_BAR(
        \g[1][11] ) );
  PG_BLOCK_594 Block_Stage_TWO_6 ( .P_ik(\p[1][13] ), .G_ik(\g[1][13] ), 
        .P_k1j(\p[1][12] ), .G_k1j(\g[1][12] ), .P_ij(\p[2][6] ), .G_ij(
        \g[2][6] ) );
  PG_BLOCK_584 Block_Stage_THREE_1 ( .P_ik(1'b0), .P_k1j(1'b0), .G_k1j(1'b0), 
        .G_ij_BAR(\g[3][1] ), .G_ik_BAR(\g[2][3] ) );
  PG_BLOCK_583 Block_Stage_THREE_2 ( .P_ik(\p[2][5] ), .G_ik(\g[2][5] ), 
        .P_k1j(\p[2][4] ), .G_k1j(\g[2][4] ), .P_ij(\p[3][2] ), .G_ij(
        \g[3][2] ) );
  G_BLOCK_166 g_4_c12_c16_1 ( .P_ik(1'b0), .G_k1j(1'b0), .G_ij(Cout[4]), 
        .G_ik_BAR(\g[3][1] ) );
  PG_BLOCK_577 Block_stage_FOUR_2_0 ( .P_ik(\p[2][6] ), .G_ik(\g[2][6] ), 
        .P_k1j(\p[3][2] ), .G_k1j(\g[3][2] ), .P_ij(\p[4][2] ), .G_ij(
        \g[4][2] ) );
  G_BLOCK_165 Block_stage_FIVE_4 ( .P_ik(\p[2][4] ), .G_ik(\g[2][4] ), .G_k1j(
        Cout[4]), .G_ij(Cout[5]) );
  G_BLOCK_164 Block_stage_FIVE_5 ( .P_ik(\p[3][2] ), .G_ik(\g[3][2] ), .G_k1j(
        Cout[4]), .G_ij(Cout[6]) );
  G_BLOCK_163 Block_stage_FIVE_6 ( .P_ik(\p[4][2] ), .G_ik(\g[4][2] ), .G_k1j(
        Cout[4]), .G_ij(Cout[7]) );
endmodule


module FA_1280 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1279 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1278 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1277 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_320 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_1280 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_1279 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_1278 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_1277 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_160 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_160 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_320 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0)
         );
  MUX_2to1_N4_160 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_1272 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1271 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1270 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1269 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_318 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_1272 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_1271 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_1270 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_1269 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_159 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_159 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_318 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0)
         );
  MUX_2to1_N4_159 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_1264 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1263 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1262 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1261 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_316 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_1264 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_1263 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_1262 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_1261 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_158 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_158 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_316 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0)
         );
  MUX_2to1_N4_158 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_1256 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1255 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1254 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1253 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_314 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1256 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1255 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1254 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1253 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_157 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_157 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_314 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  MUX_2to1_N4_157 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_1248 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1247 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1246 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1245 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_312 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1248 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1247 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1246 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1245 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1244 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_1243 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4;

  OR2_X1 U1 ( .A1(B), .A2(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(Ci), .B(n4), .ZN(S) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n4) );
  NAND2_X1 U4 ( .A1(n2), .A2(n1), .ZN(Co) );
  NAND2_X1 U5 ( .A1(B), .A2(A), .ZN(n1) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n3), .ZN(n2) );
endmodule


module FA_1242 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1241 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_311 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1244 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1243 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1242 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1241 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_156 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U3 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U4 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
endmodule


module carry_select_block_N4_156 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_312 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_311 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_156 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_1240 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1239 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1238 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4;

  OAI21_X1 U1 ( .B1(A), .B2(B), .A(Ci), .ZN(n1) );
  OAI21_X1 U2 ( .B1(n2), .B2(n3), .A(n1), .ZN(Co) );
  INV_X1 U3 ( .A(B), .ZN(n2) );
  INV_X1 U4 ( .A(A), .ZN(n3) );
  XNOR2_X1 U5 ( .A(B), .B(A), .ZN(n4) );
  XNOR2_X1 U6 ( .A(Ci), .B(n4), .ZN(S) );
endmodule


module FA_1237 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_310 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1240 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1239 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1238 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1237 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1236 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_1235 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4;

  OR2_X1 U1 ( .A1(B), .A2(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(Ci), .B(n4), .ZN(S) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n4) );
  NAND2_X1 U4 ( .A1(n2), .A2(n1), .ZN(Co) );
  NAND2_X1 U5 ( .A1(B), .A2(A), .ZN(n1) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n3), .ZN(n2) );
endmodule


module FA_1234 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1233 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(n1), .B(Ci), .ZN(S) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n1) );
endmodule


module RCA_N4_309 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1236 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1235 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1234 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1233 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_155 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
  MUX2_X2 U2 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X2 U3 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U4 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
endmodule


module carry_select_block_N4_155 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_310 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_309 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_155 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_1232 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1231 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1230 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1229 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_308 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1232 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1231 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1230 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1229 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1228 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_1227 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1226 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1225 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_307 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1228 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1227 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1226 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1225 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_154 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U3 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
  MUX2_X1 U4 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
endmodule


module carry_select_block_N4_154 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_308 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_307 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_154 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_1224 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1223 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1222 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1221 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_306 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1224 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1223 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1222 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1221 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1220 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_1219 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1218 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1217 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_305 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1220 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1219 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1218 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1217 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_153 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U3 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U4 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
endmodule


module carry_select_block_N4_153 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_306 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_305 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_153 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module SUMGENERATOR_Nblocks16_bits_per_block4_10 ( A, B, CARRY_SELECT, SUM );
  input [63:0] A;
  input [63:0] B;
  input [15:0] CARRY_SELECT;
  output [63:0] SUM;


  carry_select_block_N4_160 block_n_1 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(
        B[3:0]), .S(SUM[3:0]), .Ci(1'b0) );
  carry_select_block_N4_159 block_n_2 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(
        B[7:4]), .S(SUM[7:4]), .Ci(1'b0) );
  carry_select_block_N4_158 block_n_3 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(
        B[11:8]), .S(SUM[11:8]), .Ci(1'b0) );
  carry_select_block_N4_157 block_n_4 ( .A(A[15:12]), .B(B[15:12]), .S(
        SUM[15:12]), .Ci(1'b0) );
  carry_select_block_N4_156 block_n_5 ( .A(A[19:16]), .B(B[19:16]), .S(
        SUM[19:16]), .Ci(CARRY_SELECT[4]) );
  carry_select_block_N4_155 block_n_6 ( .A(A[23:20]), .B(B[23:20]), .S(
        SUM[23:20]), .Ci(CARRY_SELECT[5]) );
  carry_select_block_N4_154 block_n_7 ( .A(A[27:24]), .B(B[27:24]), .S(
        SUM[27:24]), .Ci(CARRY_SELECT[6]) );
  carry_select_block_N4_153 block_n_8 ( .A(A[31:28]), .B(B[31:28]), .S(
        SUM[31:28]), .Ci(CARRY_SELECT[7]) );
endmodule


module ADDER_P4_N_BIT64_10 ( A, B, add_sub, Cout, SUM );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input add_sub;
  output Cout;

  wire   [63:0] B_xor;
  wire   [15:0] tmp_co;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44;
  assign B_xor[31] = B[31];
  assign B_xor[30] = B[30];
  assign B_xor[29] = B[29];
  assign B_xor[28] = B[28];
  assign B_xor[27] = B[27];
  assign B_xor[26] = B[26];
  assign B_xor[25] = B[25];
  assign B_xor[24] = B[24];
  assign B_xor[23] = B[23];
  assign B_xor[22] = B[22];
  assign B_xor[21] = B[21];
  assign B_xor[19] = B[19];
  assign B_xor[18] = B[18];
  assign B_xor[17] = B[17];
  assign B_xor[16] = B[16];
  assign B_xor[15] = B[15];
  assign B_xor[14] = B[14];
  assign B_xor[13] = B[13];
  assign B_xor[12] = B[12];
  assign B_xor[11] = B[11];
  assign B_xor[10] = B[10];
  assign B_xor[9] = B[9];
  assign B_xor[8] = B[8];
  assign B_xor[7] = B[7];
  assign B_xor[6] = B[6];
  assign B_xor[5] = B[5];
  assign B_xor[4] = B[4];
  assign B_xor[3] = B[3];
  assign B_xor[2] = B[2];
  assign B_xor[1] = B[1];
  assign B_xor[0] = B[0];

  CARRY_GENERATOR_Nbit64_10 CLA_SPARSE_TREE ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, A[27:12], 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        B_xor[27:21], B[20], B_xor[19:12], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Cin(1'b0), .Cout({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, tmp_co[7:4], SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12}) );
  SUMGENERATOR_Nblocks16_bits_per_block4_10 CSA ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, A[31:12], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, B_xor[31:21], B[20], B_xor[19:0]}), .CARRY_SELECT({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, tmp_co[7:4], 1'b0, 
        1'b0, 1'b0, 1'b0}), .SUM({SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SUM[31:0]}) );
endmodule


module PG_NETWORK_562 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_561 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_560 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_559 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_558 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_557 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_556 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_555 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_554 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_553 ( op1, op2, g, p );
  input op1, op2;
  output g, p;
  wire   n1;

  XNOR2_X1 U1 ( .A(op2), .B(n1), .ZN(p) );
  INV_X1 U2 ( .A(op1), .ZN(n1) );
  AND2_X1 U3 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_552 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_551 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  XOR2_X1 U1 ( .A(op1), .B(op2), .Z(p) );
  AND2_X1 U2 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_550 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_549 ( op1, op2, g, p );
  input op1, op2;
  output g, p;
  wire   n1;

  INV_X1 U1 ( .A(op1), .ZN(n1) );
  XNOR2_X1 U2 ( .A(op2), .B(n1), .ZN(p) );
  AND2_X1 U3 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_BLOCK_561 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij_BAR );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij_BAR;


  AOI21_X1 U1 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(G_ij_BAR) );
endmodule


module PG_BLOCK_560 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_559 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1, n2, n3;

  INV_X1 U1 ( .A(G_ik), .ZN(n1) );
  INV_X1 U2 ( .A(P_ik), .ZN(n2) );
  INV_X1 U3 ( .A(G_k1j), .ZN(n3) );
  OAI21_X1 U4 ( .B1(n3), .B2(n2), .A(n1), .ZN(G_ij) );
  AND2_X1 U5 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
endmodule


module PG_BLOCK_558 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_557 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1, n2, n3;

  INV_X1 U1 ( .A(G_ik), .ZN(n1) );
  INV_X1 U2 ( .A(G_k1j), .ZN(n2) );
  INV_X1 U3 ( .A(P_ik), .ZN(n3) );
  OAI21_X1 U4 ( .B1(n3), .B2(n2), .A(n1), .ZN(G_ij) );
  AND2_X1 U5 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
endmodule


module PG_BLOCK_556 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(G_k1j), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_555 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1, n2;

  NAND2_X1 U1 ( .A1(n2), .A2(n1), .ZN(G_ij) );
  INV_X1 U2 ( .A(G_ik), .ZN(n1) );
  NAND2_X1 U3 ( .A1(P_ik), .A2(G_k1j), .ZN(n2) );
  AND2_X1 U4 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
endmodule


module PG_BLOCK_534 ( P_ik, P_k1j, G_k1j, P_ij, G_ij_BAR, G_ik_BAR );
  input P_ik, P_k1j, G_k1j, G_ik_BAR;
  output P_ij, G_ij_BAR;
  wire   G_ik;
  assign G_ij_BAR = G_ik;
  assign G_ik = G_ik_BAR;

endmodule


module PG_BLOCK_533 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_532 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_531 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_521 ( P_ik, P_k1j, G_k1j, P_ij, G_ij_BAR, G_ik_BAR );
  input P_ik, P_k1j, G_k1j, G_ik_BAR;
  output P_ij, G_ij_BAR;
  wire   G_ik;
  assign G_ij_BAR = G_ik;
  assign G_ik = G_ik_BAR;

endmodule


module PG_BLOCK_520 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(G_k1j), .ZN(n1) );
  OR2_X1 U2 ( .A1(G_ik), .A2(n1), .ZN(G_ij) );
  AND2_X1 U3 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
endmodule


module G_BLOCK_149 ( P_ik, G_k1j, G_ij, G_ik_BAR );
  input P_ik, G_k1j, G_ik_BAR;
  output G_ij;
  wire   G_ik;
  assign G_ik = G_ik_BAR;

  INV_X1 U1 ( .A(G_ik), .ZN(G_ij) );
endmodule


module PG_BLOCK_514 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module G_BLOCK_148 ( P_ik, G_ik, G_k1j, G_ij );
  input P_ik, G_ik, G_k1j;
  output G_ij;
  wire   n1;

  INV_X1 U1 ( .A(n1), .ZN(G_ij) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(G_k1j), .A(G_ik), .ZN(n1) );
endmodule


module G_BLOCK_147 ( P_ik, G_ik, G_k1j, G_ij );
  input P_ik, G_ik, G_k1j;
  output G_ij;
  wire   n2;

  OR2_X1 U1 ( .A1(G_ik), .A2(n2), .ZN(G_ij) );
  AND2_X1 U2 ( .A1(P_ik), .A2(G_k1j), .ZN(n2) );
endmodule


module G_BLOCK_146 ( P_ik, G_ik, G_k1j, G_ij );
  input P_ik, G_ik, G_k1j;
  output G_ij;
  wire   n1;

  OR2_X2 U1 ( .A1(G_ik), .A2(n1), .ZN(G_ij) );
  AND2_X1 U2 ( .A1(P_ik), .A2(G_k1j), .ZN(n1) );
endmodule


module CARRY_GENERATOR_Nbit64_9 ( A, B, Cin, Cout );
  input [63:0] A;
  input [63:0] B;
  output [16:0] Cout;
  input Cin;
  wire   \p[4][2] , \p[3][2] , \p[2][6] , \p[2][5] , \p[2][4] , \p[1][13] ,
         \p[1][12] , \p[1][11] , \p[1][10] , \p[1][9] , \p[1][8] , \p[0][28] ,
         \p[0][27] , \p[0][26] , \p[0][25] , \p[0][24] , \p[0][23] ,
         \p[0][22] , \p[0][21] , \p[0][20] , \p[0][19] , \p[0][18] ,
         \p[0][17] , \p[0][16] , \g[4][2] , \g[3][2] , \g[3][1] , \g[2][6] ,
         \g[2][5] , \g[2][4] , \g[2][3] , \g[1][13] , \g[1][12] , \g[1][11] ,
         \g[1][10] , \g[1][9] , \g[1][8] , \g[1][7] , \g[0][28] , \g[0][27] ,
         \g[0][26] , \g[0][25] , \g[0][24] , \g[0][23] , \g[0][22] ,
         \g[0][21] , \g[0][20] , \g[0][19] , \g[0][18] , \g[0][17] ,
         \g[0][16] , \g[0][15] ;

  PG_NETWORK_562 Block_PG_NET_15 ( .op1(A[14]), .op2(B[14]), .g(\g[0][15] ) );
  PG_NETWORK_561 Block_PG_NET_16 ( .op1(A[15]), .op2(B[15]), .g(\g[0][16] ), 
        .p(\p[0][16] ) );
  PG_NETWORK_560 Block_PG_NET_17 ( .op1(A[16]), .op2(B[16]), .g(\g[0][17] ), 
        .p(\p[0][17] ) );
  PG_NETWORK_559 Block_PG_NET_18 ( .op1(A[17]), .op2(B[17]), .g(\g[0][18] ), 
        .p(\p[0][18] ) );
  PG_NETWORK_558 Block_PG_NET_19 ( .op1(A[18]), .op2(B[18]), .g(\g[0][19] ), 
        .p(\p[0][19] ) );
  PG_NETWORK_557 Block_PG_NET_20 ( .op1(A[19]), .op2(B[19]), .g(\g[0][20] ), 
        .p(\p[0][20] ) );
  PG_NETWORK_556 Block_PG_NET_21 ( .op1(A[20]), .op2(B[20]), .g(\g[0][21] ), 
        .p(\p[0][21] ) );
  PG_NETWORK_555 Block_PG_NET_22 ( .op1(A[21]), .op2(B[21]), .g(\g[0][22] ), 
        .p(\p[0][22] ) );
  PG_NETWORK_554 Block_PG_NET_23 ( .op1(A[22]), .op2(B[22]), .g(\g[0][23] ), 
        .p(\p[0][23] ) );
  PG_NETWORK_553 Block_PG_NET_24 ( .op1(A[23]), .op2(B[23]), .g(\g[0][24] ), 
        .p(\p[0][24] ) );
  PG_NETWORK_552 Block_PG_NET_25 ( .op1(A[24]), .op2(B[24]), .g(\g[0][25] ), 
        .p(\p[0][25] ) );
  PG_NETWORK_551 Block_PG_NET_26 ( .op1(A[25]), .op2(B[25]), .g(\g[0][26] ), 
        .p(\p[0][26] ) );
  PG_NETWORK_550 Block_PG_NET_27 ( .op1(A[26]), .op2(B[26]), .g(\g[0][27] ), 
        .p(\p[0][27] ) );
  PG_NETWORK_549 Block_PG_NET_28 ( .op1(A[27]), .op2(B[27]), .g(\g[0][28] ), 
        .p(\p[0][28] ) );
  PG_BLOCK_561 Block_Stage_ONE_7 ( .P_ik(\p[0][16] ), .G_ik(\g[0][16] ), 
        .P_k1j(1'b0), .G_k1j(\g[0][15] ), .G_ij_BAR(\g[1][7] ) );
  PG_BLOCK_560 Block_Stage_ONE_8 ( .P_ik(\p[0][18] ), .G_ik(\g[0][18] ), 
        .P_k1j(\p[0][17] ), .G_k1j(\g[0][17] ), .P_ij(\p[1][8] ), .G_ij(
        \g[1][8] ) );
  PG_BLOCK_559 Block_Stage_ONE_9 ( .P_ik(\p[0][20] ), .G_ik(\g[0][20] ), 
        .P_k1j(\p[0][19] ), .G_k1j(\g[0][19] ), .P_ij(\p[1][9] ), .G_ij(
        \g[1][9] ) );
  PG_BLOCK_558 Block_Stage_ONE_10 ( .P_ik(\p[0][22] ), .G_ik(\g[0][22] ), 
        .P_k1j(\p[0][21] ), .G_k1j(\g[0][21] ), .P_ij(\p[1][10] ), .G_ij(
        \g[1][10] ) );
  PG_BLOCK_557 Block_Stage_ONE_11 ( .P_ik(\p[0][24] ), .G_ik(\g[0][24] ), 
        .P_k1j(\p[0][23] ), .G_k1j(\g[0][23] ), .P_ij(\p[1][11] ), .G_ij(
        \g[1][11] ) );
  PG_BLOCK_556 Block_Stage_ONE_12 ( .P_ik(\p[0][26] ), .G_ik(\g[0][26] ), 
        .P_k1j(\p[0][25] ), .G_k1j(\g[0][25] ), .P_ij(\p[1][12] ), .G_ij(
        \g[1][12] ) );
  PG_BLOCK_555 Block_Stage_ONE_13 ( .P_ik(\p[0][28] ), .G_ik(\g[0][28] ), 
        .P_k1j(\p[0][27] ), .G_k1j(\g[0][27] ), .P_ij(\p[1][13] ), .G_ij(
        \g[1][13] ) );
  PG_BLOCK_534 Block_Stage_TWO_3 ( .P_ik(1'b0), .P_k1j(1'b0), .G_k1j(1'b0), 
        .G_ij_BAR(\g[2][3] ), .G_ik_BAR(\g[1][7] ) );
  PG_BLOCK_533 Block_Stage_TWO_4 ( .P_ik(\p[1][9] ), .G_ik(\g[1][9] ), .P_k1j(
        \p[1][8] ), .G_k1j(\g[1][8] ), .P_ij(\p[2][4] ), .G_ij(\g[2][4] ) );
  PG_BLOCK_532 Block_Stage_TWO_5 ( .P_ik(\p[1][11] ), .G_ik(\g[1][11] ), 
        .P_k1j(\p[1][10] ), .G_k1j(\g[1][10] ), .P_ij(\p[2][5] ), .G_ij(
        \g[2][5] ) );
  PG_BLOCK_531 Block_Stage_TWO_6 ( .P_ik(\p[1][13] ), .G_ik(\g[1][13] ), 
        .P_k1j(\p[1][12] ), .G_k1j(\g[1][12] ), .P_ij(\p[2][6] ), .G_ij(
        \g[2][6] ) );
  PG_BLOCK_521 Block_Stage_THREE_1 ( .P_ik(1'b0), .P_k1j(1'b0), .G_k1j(1'b0), 
        .G_ij_BAR(\g[3][1] ), .G_ik_BAR(\g[2][3] ) );
  PG_BLOCK_520 Block_Stage_THREE_2 ( .P_ik(\p[2][5] ), .G_ik(\g[2][5] ), 
        .P_k1j(\p[2][4] ), .G_k1j(\g[2][4] ), .P_ij(\p[3][2] ), .G_ij(
        \g[3][2] ) );
  G_BLOCK_149 g_4_c12_c16_1 ( .P_ik(1'b0), .G_k1j(1'b0), .G_ij(Cout[4]), 
        .G_ik_BAR(\g[3][1] ) );
  PG_BLOCK_514 Block_stage_FOUR_2_0 ( .P_ik(\p[2][6] ), .G_ik(\g[2][6] ), 
        .P_k1j(\p[3][2] ), .G_k1j(\g[3][2] ), .P_ij(\p[4][2] ), .G_ij(
        \g[4][2] ) );
  G_BLOCK_148 Block_stage_FIVE_4 ( .P_ik(\p[2][4] ), .G_ik(\g[2][4] ), .G_k1j(
        Cout[4]), .G_ij(Cout[5]) );
  G_BLOCK_147 Block_stage_FIVE_5 ( .P_ik(\p[3][2] ), .G_ik(\g[3][2] ), .G_k1j(
        Cout[4]), .G_ij(Cout[6]) );
  G_BLOCK_146 Block_stage_FIVE_6 ( .P_ik(\p[4][2] ), .G_ik(\g[4][2] ), .G_k1j(
        Cout[4]), .G_ij(Cout[7]) );
endmodule


module FA_1152 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1151 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1150 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1149 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_288 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_1152 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_1151 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_1150 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_1149 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_144 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_144 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_288 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0)
         );
  MUX_2to1_N4_144 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_1144 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1143 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1142 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1141 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_286 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_1144 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_1143 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_1142 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_1141 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_143 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_143 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_286 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0)
         );
  MUX_2to1_N4_143 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_1136 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1135 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1134 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1133 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_284 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_1136 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_1135 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_1134 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_1133 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_142 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_142 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_284 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0)
         );
  MUX_2to1_N4_142 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_1128 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1127 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1126 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1125 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_282 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \CTMP[3] ;

  FA_1128 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_1127 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_1126 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(1'b0), .S(S[2]), .Co(\CTMP[3] ) );
  FA_1125 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(\CTMP[3] ), .S(S[3]) );
endmodule


module MUX_2to1_N4_141 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_141 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_282 RCA_0 ( .A({A[3:2], 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0) );
  MUX_2to1_N4_141 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_1120 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1119 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1118 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1117 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_280 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1120 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1119 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1118 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1117 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1116 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_1115 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1114 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1113 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_279 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1116 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1115 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1114 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1113 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_140 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U3 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U4 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
endmodule


module carry_select_block_N4_140 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_280 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_279 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_140 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_1112 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1111 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1110 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1109 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_278 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1112 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1111 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1110 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1109 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1108 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_1107 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n6) );
  XNOR2_X1 U2 ( .A(Ci), .B(n6), .ZN(S) );
  NAND2_X1 U3 ( .A1(n2), .A2(n1), .ZN(Co) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n1) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n3), .ZN(n2) );
  NAND2_X1 U6 ( .A1(n5), .A2(n4), .ZN(n3) );
  INV_X1 U7 ( .A(A), .ZN(n4) );
  INV_X1 U8 ( .A(B), .ZN(n5) );
endmodule


module FA_1106 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1105 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_277 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1108 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1107 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1106 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1105 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_139 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X2 U1 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
  MUX2_X1 U2 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U3 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U4 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
endmodule


module carry_select_block_N4_139 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_278 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_277 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_139 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_1104 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1103 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1102 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1101 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_276 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1104 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1103 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1102 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1101 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1100 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_1099 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1098 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1097 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_275 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1100 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1099 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1098 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1097 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_138 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
  MUX2_X1 U2 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U3 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U4 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
endmodule


module carry_select_block_N4_138 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_276 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_275 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_138 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_1096 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1095 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1094 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1093 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_274 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1096 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_1095 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1094 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1093 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_1092 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_1091 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1090 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_1089 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_273 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1092 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_1091 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(
        CTMP[2]) );
  FA_1090 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(
        CTMP[3]) );
  FA_1089 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_137 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X2 U1 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U3 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U4 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
endmodule


module carry_select_block_N4_137 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_274 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_273 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_137 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module SUMGENERATOR_Nblocks16_bits_per_block4_9 ( A, B, CARRY_SELECT, SUM );
  input [63:0] A;
  input [63:0] B;
  input [15:0] CARRY_SELECT;
  output [63:0] SUM;


  carry_select_block_N4_144 block_n_1 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(
        B[3:0]), .S(SUM[3:0]), .Ci(1'b0) );
  carry_select_block_N4_143 block_n_2 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(
        B[7:4]), .S(SUM[7:4]), .Ci(1'b0) );
  carry_select_block_N4_142 block_n_3 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(
        B[11:8]), .S(SUM[11:8]), .Ci(1'b0) );
  carry_select_block_N4_141 block_n_4 ( .A({A[15:14], 1'b0, 1'b0}), .B(
        B[15:12]), .S(SUM[15:12]), .Ci(1'b0) );
  carry_select_block_N4_140 block_n_5 ( .A(A[19:16]), .B(B[19:16]), .S(
        SUM[19:16]), .Ci(CARRY_SELECT[4]) );
  carry_select_block_N4_139 block_n_6 ( .A(A[23:20]), .B(B[23:20]), .S(
        SUM[23:20]), .Ci(CARRY_SELECT[5]) );
  carry_select_block_N4_138 block_n_7 ( .A(A[27:24]), .B(B[27:24]), .S(
        SUM[27:24]), .Ci(CARRY_SELECT[6]) );
  carry_select_block_N4_137 block_n_8 ( .A(A[31:28]), .B(B[31:28]), .S(
        SUM[31:28]), .Ci(CARRY_SELECT[7]) );
endmodule


module ADDER_P4_N_BIT64_9 ( A, B, add_sub, Cout, SUM );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input add_sub;
  output Cout;
  wire   n1;
  wire   [63:0] B_xor;
  wire   [15:0] tmp_co;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44;
  assign B_xor[31] = B[31];
  assign B_xor[30] = B[30];
  assign B_xor[29] = B[29];
  assign B_xor[28] = B[28];
  assign B_xor[27] = B[27];
  assign B_xor[26] = B[26];
  assign B_xor[25] = B[25];
  assign B_xor[24] = B[24];
  assign B_xor[23] = B[23];
  assign B_xor[22] = B[22];
  assign B_xor[21] = B[21];
  assign B_xor[20] = B[20];
  assign B_xor[19] = B[19];
  assign B_xor[18] = B[18];
  assign B_xor[17] = B[17];
  assign B_xor[16] = B[16];
  assign B_xor[15] = B[15];
  assign B_xor[14] = B[14];
  assign B_xor[13] = B[13];
  assign B_xor[12] = B[12];
  assign B_xor[11] = B[11];
  assign B_xor[10] = B[10];
  assign B_xor[9] = B[9];
  assign B_xor[8] = B[8];
  assign B_xor[7] = B[7];
  assign B_xor[6] = B[6];
  assign B_xor[5] = B[5];
  assign B_xor[4] = B[4];
  assign B_xor[3] = B[3];
  assign B_xor[2] = B[2];
  assign B_xor[1] = B[1];
  assign B_xor[0] = B[0];

  CARRY_GENERATOR_Nbit64_9 CLA_SPARSE_TREE ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, A[27:14], 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, B_xor[27:14], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Cin(1'b0), .Cout({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, tmp_co[7:4], SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12}) );
  SUMGENERATOR_Nblocks16_bits_per_block4_9 CSA ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, A[31:14], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B_xor[31:26], n1, B_xor[24:0]}), 
        .CARRY_SELECT({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        tmp_co[7:4], 1'b0, 1'b0, 1'b0, 1'b0}), .SUM({SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SUM[31:0]}) );
  BUF_X1 U1 ( .A(B_xor[25]), .Z(n1) );
endmodule


module PG_NETWORK_496 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_495 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_494 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_493 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_492 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_491 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_490 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_489 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_488 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_487 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  XOR2_X1 U1 ( .A(op1), .B(op2), .Z(p) );
  AND2_X1 U2 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_486 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_485 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  XOR2_X1 U1 ( .A(op1), .B(op2), .Z(p) );
  AND2_X1 U2 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_BLOCK_497 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AOI21_X1 U1 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_496 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_495 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_494 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_493 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_492 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij_BAR );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij_BAR;


  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(G_k1j), .A(G_ik), .ZN(G_ij_BAR) );
endmodule


module PG_BLOCK_470 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij_BAR );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij_BAR;


  AOI21_X1 U1 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(G_ij_BAR) );
endmodule


module PG_BLOCK_469 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_468 ( P_ik, P_k1j, G_k1j, P_ij, G_ij, G_ik_BAR );
  input P_ik, P_k1j, G_k1j, G_ik_BAR;
  output P_ij, G_ij;
  wire   G_ik, n1;
  assign G_ik = G_ik_BAR;

  NAND2_X1 U1 ( .A1(n1), .A2(G_ik), .ZN(G_ij) );
  NAND2_X1 U2 ( .A1(G_k1j), .A2(P_ik), .ZN(n1) );
  AND2_X1 U3 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
endmodule


module PG_BLOCK_457 ( P_ik, G_ik, P_k1j, P_ij, G_ij_BAR, G_k1j_BAR );
  input P_ik, G_ik, P_k1j, G_k1j_BAR;
  output P_ij, G_ij_BAR;
  wire   G_k1j, n1;
  assign G_k1j = G_k1j_BAR;

  INV_X1 U1 ( .A(G_k1j), .ZN(n1) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(n1), .A(G_ik), .ZN(G_ij_BAR) );
endmodule


module PG_BLOCK_451 ( P_ik, G_ik, P_k1j, P_ij, G_ij_BAR, G_k1j_BAR );
  input P_ik, G_ik, P_k1j, G_k1j_BAR;
  output P_ij, G_ij_BAR;
  wire   G_k1j, n1;
  assign G_k1j = G_k1j_BAR;

  INV_X1 U1 ( .A(G_k1j), .ZN(n1) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(n1), .A(G_ik), .ZN(G_ij_BAR) );
endmodule


module G_BLOCK_131 ( P_ik, G_k1j, G_ij, G_ik_BAR );
  input P_ik, G_k1j, G_ik_BAR;
  output G_ij;
  wire   G_ik;
  assign G_ik = G_ik_BAR;

  INV_X1 U1 ( .A(G_ik), .ZN(G_ij) );
endmodule


module G_BLOCK_130 ( P_ik, G_k1j, G_ij, G_ik_BAR );
  input P_ik, G_k1j, G_ik_BAR;
  output G_ij;
  wire   G_ik;
  assign G_ik = G_ik_BAR;

  INV_X1 U1 ( .A(G_ik), .ZN(G_ij) );
endmodule


module G_BLOCK_129 ( P_ik, G_k1j, G_ij, G_ik_BAR );
  input P_ik, G_k1j, G_ik_BAR;
  output G_ij;
  wire   G_ik;
  assign G_ik = G_ik_BAR;

  INV_X1 U1 ( .A(G_ik), .ZN(G_ij) );
endmodule


module CARRY_GENERATOR_Nbit64_8 ( A, B, Cin, Cout );
  input [63:0] A;
  input [63:0] B;
  output [16:0] Cout;
  input Cin;
  wire   \p[2][6] , \p[2][5] , \p[1][13] , \p[1][12] , \p[1][11] , \p[1][10] ,
         \p[1][9] , \p[0][28] , \p[0][27] , \p[0][26] , \p[0][25] , \p[0][24] ,
         \p[0][23] , \p[0][22] , \p[0][21] , \p[0][20] , \p[0][19] ,
         \p[0][18] , \g[4][2] , \g[3][2] , \g[2][6] , \g[2][5] , \g[2][4] ,
         \g[1][13] , \g[1][12] , \g[1][11] , \g[1][10] , \g[1][9] , \g[1][8] ,
         \g[0][28] , \g[0][27] , \g[0][26] , \g[0][25] , \g[0][24] ,
         \g[0][23] , \g[0][22] , \g[0][21] , \g[0][20] , \g[0][19] ,
         \g[0][18] , \g[0][17] , n1;

  PG_NETWORK_496 Block_PG_NET_17 ( .op1(A[16]), .op2(B[16]), .g(\g[0][17] ) );
  PG_NETWORK_495 Block_PG_NET_18 ( .op1(A[17]), .op2(B[17]), .g(\g[0][18] ), 
        .p(\p[0][18] ) );
  PG_NETWORK_494 Block_PG_NET_19 ( .op1(A[18]), .op2(B[18]), .g(\g[0][19] ), 
        .p(\p[0][19] ) );
  PG_NETWORK_493 Block_PG_NET_20 ( .op1(A[19]), .op2(B[19]), .g(\g[0][20] ), 
        .p(\p[0][20] ) );
  PG_NETWORK_492 Block_PG_NET_21 ( .op1(A[20]), .op2(B[20]), .g(\g[0][21] ), 
        .p(\p[0][21] ) );
  PG_NETWORK_491 Block_PG_NET_22 ( .op1(A[21]), .op2(B[21]), .g(\g[0][22] ), 
        .p(\p[0][22] ) );
  PG_NETWORK_490 Block_PG_NET_23 ( .op1(A[22]), .op2(B[22]), .g(\g[0][23] ), 
        .p(\p[0][23] ) );
  PG_NETWORK_489 Block_PG_NET_24 ( .op1(A[23]), .op2(B[23]), .g(\g[0][24] ), 
        .p(\p[0][24] ) );
  PG_NETWORK_488 Block_PG_NET_25 ( .op1(A[24]), .op2(B[24]), .g(\g[0][25] ), 
        .p(\p[0][25] ) );
  PG_NETWORK_487 Block_PG_NET_26 ( .op1(A[25]), .op2(B[25]), .g(\g[0][26] ), 
        .p(\p[0][26] ) );
  PG_NETWORK_486 Block_PG_NET_27 ( .op1(A[26]), .op2(B[26]), .g(\g[0][27] ), 
        .p(\p[0][27] ) );
  PG_NETWORK_485 Block_PG_NET_28 ( .op1(A[27]), .op2(B[27]), .g(\g[0][28] ), 
        .p(\p[0][28] ) );
  PG_BLOCK_497 Block_Stage_ONE_8 ( .P_ik(\p[0][18] ), .G_ik(\g[0][18] ), 
        .P_k1j(1'b0), .G_k1j(\g[0][17] ), .G_ij(\g[1][8] ) );
  PG_BLOCK_496 Block_Stage_ONE_9 ( .P_ik(\p[0][20] ), .G_ik(\g[0][20] ), 
        .P_k1j(\p[0][19] ), .G_k1j(\g[0][19] ), .P_ij(\p[1][9] ), .G_ij(
        \g[1][9] ) );
  PG_BLOCK_495 Block_Stage_ONE_10 ( .P_ik(\p[0][22] ), .G_ik(\g[0][22] ), 
        .P_k1j(\p[0][21] ), .G_k1j(\g[0][21] ), .P_ij(\p[1][10] ), .G_ij(
        \g[1][10] ) );
  PG_BLOCK_494 Block_Stage_ONE_11 ( .P_ik(\p[0][24] ), .G_ik(\g[0][24] ), 
        .P_k1j(\p[0][23] ), .G_k1j(\g[0][23] ), .P_ij(\p[1][11] ), .G_ij(
        \g[1][11] ) );
  PG_BLOCK_493 Block_Stage_ONE_12 ( .P_ik(\p[0][26] ), .G_ik(\g[0][26] ), 
        .P_k1j(\p[0][25] ), .G_k1j(\g[0][25] ), .P_ij(\p[1][12] ), .G_ij(
        \g[1][12] ) );
  PG_BLOCK_492 Block_Stage_ONE_13 ( .P_ik(\p[0][28] ), .G_ik(\g[0][28] ), 
        .P_k1j(\p[0][27] ), .G_k1j(\g[0][27] ), .P_ij(\p[1][13] ), .G_ij_BAR(
        \g[1][13] ) );
  PG_BLOCK_470 Block_Stage_TWO_4 ( .P_ik(\p[1][9] ), .G_ik(\g[1][9] ), .P_k1j(
        1'b0), .G_k1j(\g[1][8] ), .G_ij_BAR(\g[2][4] ) );
  PG_BLOCK_469 Block_Stage_TWO_5 ( .P_ik(\p[1][11] ), .G_ik(\g[1][11] ), 
        .P_k1j(\p[1][10] ), .G_k1j(\g[1][10] ), .P_ij(\p[2][5] ), .G_ij(
        \g[2][5] ) );
  PG_BLOCK_468 Block_Stage_TWO_6 ( .P_ik(\p[1][13] ), .P_k1j(\p[1][12] ), 
        .G_k1j(\g[1][12] ), .P_ij(\p[2][6] ), .G_ij(\g[2][6] ), .G_ik_BAR(
        \g[1][13] ) );
  PG_BLOCK_457 Block_Stage_THREE_2 ( .P_ik(\p[2][5] ), .G_ik(\g[2][5] ), 
        .P_k1j(1'b0), .G_ij_BAR(\g[3][2] ), .G_k1j_BAR(\g[2][4] ) );
  PG_BLOCK_451 Block_stage_FOUR_2_0 ( .P_ik(\p[2][6] ), .G_ik(\g[2][6] ), 
        .P_k1j(1'b0), .G_ij_BAR(\g[4][2] ), .G_k1j_BAR(\g[3][2] ) );
  G_BLOCK_131 Block_stage_FIVE_4 ( .P_ik(1'b0), .G_k1j(1'b0), .G_ij(Cout[5]), 
        .G_ik_BAR(\g[2][4] ) );
  G_BLOCK_130 Block_stage_FIVE_5 ( .P_ik(1'b0), .G_k1j(1'b0), .G_ij(Cout[6]), 
        .G_ik_BAR(n1) );
  G_BLOCK_129 Block_stage_FIVE_6 ( .P_ik(1'b0), .G_k1j(1'b0), .G_ij(Cout[7]), 
        .G_ik_BAR(\g[4][2] ) );
  BUF_X1 U1 ( .A(\g[3][2] ), .Z(n1) );
endmodule


module FA_1024 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1023 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1022 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1021 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_256 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_1024 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_1023 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_1022 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_1021 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_128 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_128 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_256 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0)
         );
  MUX_2to1_N4_128 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_1016 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1015 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1014 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1013 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_254 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_1016 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_1015 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_1014 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_1013 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_127 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_127 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_254 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0)
         );
  MUX_2to1_N4_127 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_1008 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1007 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1006 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_1005 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_252 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_1008 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_1007 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_1006 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_1005 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_126 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_126 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_252 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0)
         );
  MUX_2to1_N4_126 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_1000 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_999 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_998 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_997 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_250 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_1000 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_999 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_998 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_997 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_125 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_125 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_250 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0)
         );
  MUX_2to1_N4_125 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_992 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_991 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_990 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_989 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_248 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_992 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_991 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_990 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_989 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_124 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_124 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_248 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  MUX_2to1_N4_124 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_984 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_983 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_982 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_981 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_246 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_984 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_983 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_982 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_981 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_980 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_979 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_978 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_977 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_245 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_980 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_979 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_978 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_977 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_123 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U3 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U4 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
endmodule


module carry_select_block_N4_123 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_246 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_245 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_123 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_976 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_975 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_974 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_973 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_244 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_976 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_975 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_974 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_973 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_972 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_971 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_970 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_969 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_243 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_972 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_971 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_970 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_969 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_122 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;
  wire   n1, n2, n3;

  NAND2_X1 U1 ( .A1(n3), .A2(n1), .ZN(Y[3]) );
  NAND2_X1 U2 ( .A1(IN0[3]), .A2(n2), .ZN(n1) );
  INV_X1 U3 ( .A(SEL), .ZN(n2) );
  NAND2_X1 U4 ( .A1(IN1[3]), .A2(SEL), .ZN(n3) );
  MUX2_X1 U5 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U6 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U7 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
endmodule


module carry_select_block_N4_122 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_244 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_243 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_122 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_968 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_967 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_966 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4;

  OR2_X1 U1 ( .A1(B), .A2(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(Ci), .B(n4), .ZN(S) );
  NAND2_X1 U3 ( .A1(n2), .A2(n1), .ZN(Co) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n2) );
  NAND2_X1 U5 ( .A1(B), .A2(A), .ZN(n1) );
  XNOR2_X1 U6 ( .A(B), .B(A), .ZN(n4) );
endmodule


module FA_965 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_242 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_968 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_967 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_966 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_965 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_964 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_963 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(Ci), .B(n6), .ZN(S) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(n2), .A2(n1), .ZN(Co) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n1) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n3), .ZN(n2) );
  NAND2_X1 U6 ( .A1(n5), .A2(n4), .ZN(n3) );
  INV_X1 U7 ( .A(A), .ZN(n4) );
  INV_X1 U8 ( .A(B), .ZN(n5) );
endmodule


module FA_962 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(Ci), .B(n6), .ZN(S) );
  NAND2_X1 U2 ( .A1(n2), .A2(n1), .ZN(Co) );
  NAND2_X1 U3 ( .A1(Ci), .A2(n3), .ZN(n2) );
  NAND2_X1 U4 ( .A1(n5), .A2(n4), .ZN(n3) );
  INV_X1 U5 ( .A(B), .ZN(n5) );
  NAND2_X1 U6 ( .A1(B), .A2(A), .ZN(n1) );
  XNOR2_X1 U7 ( .A(B), .B(A), .ZN(n6) );
  INV_X1 U8 ( .A(A), .ZN(n4) );
endmodule


module FA_961 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(Ci), .B(n1), .ZN(S) );
endmodule


module RCA_N4_241 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_964 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_963 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_962 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_961 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_121 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U3 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U4 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
endmodule


module carry_select_block_N4_121 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_242 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_241 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_121 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module SUMGENERATOR_Nblocks16_bits_per_block4_8 ( A, B, CARRY_SELECT, SUM );
  input [63:0] A;
  input [63:0] B;
  input [15:0] CARRY_SELECT;
  output [63:0] SUM;


  carry_select_block_N4_128 block_n_1 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(
        B[3:0]), .S(SUM[3:0]), .Ci(1'b0) );
  carry_select_block_N4_127 block_n_2 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(
        B[7:4]), .S(SUM[7:4]), .Ci(1'b0) );
  carry_select_block_N4_126 block_n_3 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(
        B[11:8]), .S(SUM[11:8]), .Ci(1'b0) );
  carry_select_block_N4_125 block_n_4 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(
        B[15:12]), .S(SUM[15:12]), .Ci(1'b0) );
  carry_select_block_N4_124 block_n_5 ( .A(A[19:16]), .B(B[19:16]), .S(
        SUM[19:16]), .Ci(1'b0) );
  carry_select_block_N4_123 block_n_6 ( .A(A[23:20]), .B(B[23:20]), .S(
        SUM[23:20]), .Ci(CARRY_SELECT[5]) );
  carry_select_block_N4_122 block_n_7 ( .A(A[27:24]), .B(B[27:24]), .S(
        SUM[27:24]), .Ci(CARRY_SELECT[6]) );
  carry_select_block_N4_121 block_n_8 ( .A(A[31:28]), .B(B[31:28]), .S(
        SUM[31:28]), .Ci(CARRY_SELECT[7]) );
endmodule


module ADDER_P4_N_BIT64_8 ( A, B, add_sub, Cout, SUM );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input add_sub;
  output Cout;

  wire   [63:0] B_xor;
  wire   [15:0] tmp_co;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45;
  assign B_xor[31] = B[31];
  assign B_xor[30] = B[30];
  assign B_xor[29] = B[29];
  assign B_xor[27] = B[27];
  assign B_xor[26] = B[26];
  assign B_xor[25] = B[25];
  assign B_xor[24] = B[24];
  assign B_xor[23] = B[23];
  assign B_xor[22] = B[22];
  assign B_xor[21] = B[21];
  assign B_xor[20] = B[20];
  assign B_xor[19] = B[19];
  assign B_xor[18] = B[18];
  assign B_xor[17] = B[17];
  assign B_xor[16] = B[16];
  assign B_xor[15] = B[15];
  assign B_xor[14] = B[14];
  assign B_xor[13] = B[13];
  assign B_xor[12] = B[12];
  assign B_xor[11] = B[11];
  assign B_xor[10] = B[10];
  assign B_xor[9] = B[9];
  assign B_xor[8] = B[8];
  assign B_xor[7] = B[7];
  assign B_xor[6] = B[6];
  assign B_xor[5] = B[5];
  assign B_xor[4] = B[4];
  assign B_xor[3] = B[3];
  assign B_xor[2] = B[2];
  assign B_xor[1] = B[1];
  assign B_xor[0] = B[0];

  CARRY_GENERATOR_Nbit64_8 CLA_SPARSE_TREE ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, A[27:16], 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, B_xor[27:16], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Cin(1'b0), 
        .Cout({SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, tmp_co[7:5], SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13}) );
  SUMGENERATOR_Nblocks16_bits_per_block4_8 CSA ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, A[31:16], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B_xor[31:29], B[28], 
        B_xor[27:0]}), .CARRY_SELECT({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, tmp_co[7:5], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .SUM({
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, SUM[31:0]}) );
endmodule


module PG_NETWORK_430 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_429 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_428 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_427 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_426 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_425 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_424 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_423 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_422 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_421 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_BLOCK_433 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij_BAR );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij_BAR;


  AOI21_X1 U1 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(G_ij_BAR) );
endmodule


module PG_BLOCK_432 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_431 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_430 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_429 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_407 ( P_ik, P_k1j, G_k1j, P_ij, G_ij_BAR, G_ik_BAR );
  input P_ik, P_k1j, G_k1j, G_ik_BAR;
  output P_ij, G_ij_BAR;
  wire   G_ik;
  assign G_ij_BAR = G_ik;
  assign G_ik = G_ik_BAR;

endmodule


module PG_BLOCK_406 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_405 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_394 ( P_ik, G_ik, P_k1j, P_ij, G_ij_BAR, G_k1j_BAR );
  input P_ik, G_ik, P_k1j, G_k1j_BAR;
  output P_ij, G_ij_BAR;
  wire   G_k1j, n1;
  assign G_k1j = G_k1j_BAR;

  INV_X1 U1 ( .A(G_k1j), .ZN(n1) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(n1), .A(G_ik), .ZN(G_ij_BAR) );
endmodule


module PG_BLOCK_388 ( P_ik, G_ik, P_k1j, P_ij, G_ij_BAR, G_k1j_BAR );
  input P_ik, G_ik, P_k1j, G_k1j_BAR;
  output P_ij, G_ij_BAR;
  wire   G_k1j, n1;
  assign G_k1j = G_k1j_BAR;

  INV_X1 U1 ( .A(G_k1j), .ZN(n1) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(n1), .A(G_ik), .ZN(G_ij_BAR) );
endmodule


module G_BLOCK_114 ( P_ik, G_k1j, G_ij, G_ik_BAR );
  input P_ik, G_k1j, G_ik_BAR;
  output G_ij;
  wire   G_ik;
  assign G_ik = G_ik_BAR;

  INV_X1 U1 ( .A(G_ik), .ZN(G_ij) );
endmodule


module G_BLOCK_113 ( P_ik, G_k1j, G_ij, G_ik_BAR );
  input P_ik, G_k1j, G_ik_BAR;
  output G_ij;
  wire   G_ik;
  assign G_ik = G_ik_BAR;

  INV_X1 U1 ( .A(G_ik), .ZN(G_ij) );
endmodule


module G_BLOCK_112 ( P_ik, G_k1j, G_ij, G_ik_BAR );
  input P_ik, G_k1j, G_ik_BAR;
  output G_ij;
  wire   G_ik;
  assign G_ik = G_ik_BAR;

  INV_X1 U1 ( .A(G_ik), .ZN(G_ij) );
endmodule


module CARRY_GENERATOR_Nbit64_7 ( A, B, Cin, Cout );
  input [63:0] A;
  input [63:0] B;
  output [16:0] Cout;
  input Cin;
  wire   \p[2][6] , \p[2][5] , \p[1][13] , \p[1][12] , \p[1][11] , \p[1][10] ,
         \p[0][28] , \p[0][27] , \p[0][26] , \p[0][25] , \p[0][24] ,
         \p[0][23] , \p[0][22] , \p[0][21] , \p[0][20] , \g[4][2] , \g[3][2] ,
         \g[2][6] , \g[2][5] , \g[2][4] , \g[1][13] , \g[1][12] , \g[1][11] ,
         \g[1][10] , \g[1][9] , \g[0][28] , \g[0][27] , \g[0][26] , \g[0][25] ,
         \g[0][24] , \g[0][23] , \g[0][22] , \g[0][21] , \g[0][20] ,
         \g[0][19] ;

  PG_NETWORK_430 Block_PG_NET_19 ( .op1(A[18]), .op2(B[18]), .g(\g[0][19] ) );
  PG_NETWORK_429 Block_PG_NET_20 ( .op1(A[19]), .op2(B[19]), .g(\g[0][20] ), 
        .p(\p[0][20] ) );
  PG_NETWORK_428 Block_PG_NET_21 ( .op1(A[20]), .op2(B[20]), .g(\g[0][21] ), 
        .p(\p[0][21] ) );
  PG_NETWORK_427 Block_PG_NET_22 ( .op1(A[21]), .op2(B[21]), .g(\g[0][22] ), 
        .p(\p[0][22] ) );
  PG_NETWORK_426 Block_PG_NET_23 ( .op1(A[22]), .op2(B[22]), .g(\g[0][23] ), 
        .p(\p[0][23] ) );
  PG_NETWORK_425 Block_PG_NET_24 ( .op1(A[23]), .op2(B[23]), .g(\g[0][24] ), 
        .p(\p[0][24] ) );
  PG_NETWORK_424 Block_PG_NET_25 ( .op1(A[24]), .op2(B[24]), .g(\g[0][25] ), 
        .p(\p[0][25] ) );
  PG_NETWORK_423 Block_PG_NET_26 ( .op1(A[25]), .op2(B[25]), .g(\g[0][26] ), 
        .p(\p[0][26] ) );
  PG_NETWORK_422 Block_PG_NET_27 ( .op1(A[26]), .op2(B[26]), .g(\g[0][27] ), 
        .p(\p[0][27] ) );
  PG_NETWORK_421 Block_PG_NET_28 ( .op1(A[27]), .op2(B[27]), .g(\g[0][28] ), 
        .p(\p[0][28] ) );
  PG_BLOCK_433 Block_Stage_ONE_9 ( .P_ik(\p[0][20] ), .G_ik(\g[0][20] ), 
        .P_k1j(1'b0), .G_k1j(\g[0][19] ), .G_ij_BAR(\g[1][9] ) );
  PG_BLOCK_432 Block_Stage_ONE_10 ( .P_ik(\p[0][22] ), .G_ik(\g[0][22] ), 
        .P_k1j(\p[0][21] ), .G_k1j(\g[0][21] ), .P_ij(\p[1][10] ), .G_ij(
        \g[1][10] ) );
  PG_BLOCK_431 Block_Stage_ONE_11 ( .P_ik(\p[0][24] ), .G_ik(\g[0][24] ), 
        .P_k1j(\p[0][23] ), .G_k1j(\g[0][23] ), .P_ij(\p[1][11] ), .G_ij(
        \g[1][11] ) );
  PG_BLOCK_430 Block_Stage_ONE_12 ( .P_ik(\p[0][26] ), .G_ik(\g[0][26] ), 
        .P_k1j(\p[0][25] ), .G_k1j(\g[0][25] ), .P_ij(\p[1][12] ), .G_ij(
        \g[1][12] ) );
  PG_BLOCK_429 Block_Stage_ONE_13 ( .P_ik(\p[0][28] ), .G_ik(\g[0][28] ), 
        .P_k1j(\p[0][27] ), .G_k1j(\g[0][27] ), .P_ij(\p[1][13] ), .G_ij(
        \g[1][13] ) );
  PG_BLOCK_407 Block_Stage_TWO_4 ( .P_ik(1'b0), .P_k1j(1'b0), .G_k1j(1'b0), 
        .G_ij_BAR(\g[2][4] ), .G_ik_BAR(\g[1][9] ) );
  PG_BLOCK_406 Block_Stage_TWO_5 ( .P_ik(\p[1][11] ), .G_ik(\g[1][11] ), 
        .P_k1j(\p[1][10] ), .G_k1j(\g[1][10] ), .P_ij(\p[2][5] ), .G_ij(
        \g[2][5] ) );
  PG_BLOCK_405 Block_Stage_TWO_6 ( .P_ik(\p[1][13] ), .G_ik(\g[1][13] ), 
        .P_k1j(\p[1][12] ), .G_k1j(\g[1][12] ), .P_ij(\p[2][6] ), .G_ij(
        \g[2][6] ) );
  PG_BLOCK_394 Block_Stage_THREE_2 ( .P_ik(\p[2][5] ), .G_ik(\g[2][5] ), 
        .P_k1j(1'b0), .G_ij_BAR(\g[3][2] ), .G_k1j_BAR(\g[2][4] ) );
  PG_BLOCK_388 Block_stage_FOUR_2_0 ( .P_ik(\p[2][6] ), .G_ik(\g[2][6] ), 
        .P_k1j(1'b0), .G_ij_BAR(\g[4][2] ), .G_k1j_BAR(\g[3][2] ) );
  G_BLOCK_114 Block_stage_FIVE_4 ( .P_ik(1'b0), .G_k1j(1'b0), .G_ij(Cout[5]), 
        .G_ik_BAR(\g[2][4] ) );
  G_BLOCK_113 Block_stage_FIVE_5 ( .P_ik(1'b0), .G_k1j(1'b0), .G_ij(Cout[6]), 
        .G_ik_BAR(\g[3][2] ) );
  G_BLOCK_112 Block_stage_FIVE_6 ( .P_ik(1'b0), .G_k1j(1'b0), .G_ij(Cout[7]), 
        .G_ik_BAR(\g[4][2] ) );
endmodule


module FA_896 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_895 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_894 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_893 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_224 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_896 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_895 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_894 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_893 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_112 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_112 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_224 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0)
         );
  MUX_2to1_N4_112 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_888 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_887 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_886 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_885 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_222 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_888 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_887 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_886 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_885 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_111 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_111 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_222 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0)
         );
  MUX_2to1_N4_111 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_880 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_879 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_878 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_877 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_220 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_880 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_879 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_878 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_877 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_110 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_110 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_220 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0)
         );
  MUX_2to1_N4_110 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_872 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_871 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_870 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_869 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_218 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_872 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_871 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_870 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_869 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_109 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_109 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_218 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0)
         );
  MUX_2to1_N4_109 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_864 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_863 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_862 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_861 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_216 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \CTMP[3] ;

  FA_864 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_863 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_862 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(1'b0), .S(S[2]), .Co(\CTMP[3] )
         );
  FA_861 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(\CTMP[3] ), .S(S[3]) );
endmodule


module MUX_2to1_N4_108 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_108 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_216 RCA_0 ( .A({A[3:2], 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0) );
  MUX_2to1_N4_108 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_856 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_855 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_854 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_853 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_214 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_856 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_855 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_854 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_853 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_852 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_851 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_850 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_849 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_213 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_852 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_851 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_850 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_849 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_107 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U3 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U4 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
endmodule


module carry_select_block_N4_107 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_214 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_213 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_107 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_848 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_847 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_846 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_845 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_212 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_848 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_847 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_846 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_845 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_844 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_843 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_842 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_841 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_211 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_844 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_843 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_842 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_841 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_106 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U3 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U4 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
endmodule


module carry_select_block_N4_106 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_212 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_211 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_106 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_840 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_839 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_838 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_837 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_210 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_840 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_839 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_838 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_837 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_836 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_835 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_834 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_833 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_209 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_836 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_835 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_834 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_833 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_105 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U3 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U4 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
endmodule


module carry_select_block_N4_105 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_210 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_209 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_105 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module SUMGENERATOR_Nblocks16_bits_per_block4_7 ( A, B, CARRY_SELECT, SUM );
  input [63:0] A;
  input [63:0] B;
  input [15:0] CARRY_SELECT;
  output [63:0] SUM;


  carry_select_block_N4_112 block_n_1 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(
        B[3:0]), .S(SUM[3:0]), .Ci(1'b0) );
  carry_select_block_N4_111 block_n_2 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(
        B[7:4]), .S(SUM[7:4]), .Ci(1'b0) );
  carry_select_block_N4_110 block_n_3 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(
        B[11:8]), .S(SUM[11:8]), .Ci(1'b0) );
  carry_select_block_N4_109 block_n_4 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(
        B[15:12]), .S(SUM[15:12]), .Ci(1'b0) );
  carry_select_block_N4_108 block_n_5 ( .A({A[19:18], 1'b0, 1'b0}), .B(
        B[19:16]), .S(SUM[19:16]), .Ci(1'b0) );
  carry_select_block_N4_107 block_n_6 ( .A(A[23:20]), .B(B[23:20]), .S(
        SUM[23:20]), .Ci(CARRY_SELECT[5]) );
  carry_select_block_N4_106 block_n_7 ( .A(A[27:24]), .B(B[27:24]), .S(
        SUM[27:24]), .Ci(CARRY_SELECT[6]) );
  carry_select_block_N4_105 block_n_8 ( .A(A[31:28]), .B(B[31:28]), .S(
        SUM[31:28]), .Ci(CARRY_SELECT[7]) );
endmodule


module ADDER_P4_N_BIT64_7 ( A, B, add_sub, Cout, SUM );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input add_sub;
  output Cout;

  wire   [63:0] B_xor;
  wire   [15:0] tmp_co;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45;
  assign B_xor[31] = B[31];
  assign B_xor[30] = B[30];
  assign B_xor[29] = B[29];
  assign B_xor[28] = B[28];
  assign B_xor[27] = B[27];
  assign B_xor[26] = B[26];
  assign B_xor[25] = B[25];
  assign B_xor[24] = B[24];
  assign B_xor[23] = B[23];
  assign B_xor[22] = B[22];
  assign B_xor[21] = B[21];
  assign B_xor[20] = B[20];
  assign B_xor[19] = B[19];
  assign B_xor[18] = B[18];
  assign B_xor[17] = B[17];
  assign B_xor[16] = B[16];
  assign B_xor[15] = B[15];
  assign B_xor[14] = B[14];
  assign B_xor[13] = B[13];
  assign B_xor[12] = B[12];
  assign B_xor[11] = B[11];
  assign B_xor[10] = B[10];
  assign B_xor[9] = B[9];
  assign B_xor[8] = B[8];
  assign B_xor[7] = B[7];
  assign B_xor[6] = B[6];
  assign B_xor[5] = B[5];
  assign B_xor[4] = B[4];
  assign B_xor[3] = B[3];
  assign B_xor[2] = B[2];
  assign B_xor[1] = B[1];
  assign B_xor[0] = B[0];

  CARRY_GENERATOR_Nbit64_7 CLA_SPARSE_TREE ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, A[27:18], 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, B_xor[27:18], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .Cin(1'b0), .Cout({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, tmp_co[7:5], 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13}) );
  SUMGENERATOR_Nblocks16_bits_per_block4_7 CSA ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, A[31:18], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B_xor[31:0]}), 
        .CARRY_SELECT({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        tmp_co[7:5], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .SUM({
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, SUM[31:0]}) );
endmodule


module PG_NETWORK_364 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_363 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_362 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_361 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_360 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_359 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_358 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_357 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_BLOCK_369 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AOI21_X1 U1 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_368 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_367 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_366 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_343 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij_BAR );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij_BAR;


  AOI21_X1 U1 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(G_ij_BAR) );
endmodule


module PG_BLOCK_342 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_331 ( P_ik, P_k1j, G_k1j, P_ij, G_ij_BAR, G_ik_BAR );
  input P_ik, P_k1j, G_k1j, G_ik_BAR;
  output P_ij, G_ij_BAR;
  wire   G_ik;
  assign G_ij_BAR = G_ik;
  assign G_ik = G_ik_BAR;

endmodule


module PG_BLOCK_325 ( P_ik, G_ik, P_k1j, P_ij, G_ij_BAR, G_k1j_BAR );
  input P_ik, G_ik, P_k1j, G_k1j_BAR;
  output P_ij, G_ij_BAR;
  wire   G_k1j, n1;
  assign G_k1j = G_k1j_BAR;

  INV_X1 U1 ( .A(G_k1j), .ZN(n1) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(n1), .A(G_ik), .ZN(G_ij_BAR) );
endmodule


module G_BLOCK_96 ( P_ik, G_k1j, G_ij, G_ik_BAR );
  input P_ik, G_k1j, G_ik_BAR;
  output G_ij;
  wire   G_ik;
  assign G_ik = G_ik_BAR;

  INV_X1 U1 ( .A(G_ik), .ZN(G_ij) );
endmodule


module G_BLOCK_95 ( P_ik, G_k1j, G_ij, G_ik_BAR );
  input P_ik, G_k1j, G_ik_BAR;
  output G_ij;
  wire   G_ik;
  assign G_ik = G_ik_BAR;

  INV_X1 U1 ( .A(G_ik), .ZN(G_ij) );
endmodule


module CARRY_GENERATOR_Nbit64_6 ( A, B, Cin, Cout );
  input [63:0] A;
  input [63:0] B;
  output [16:0] Cout;
  input Cin;
  wire   \p[2][6] , \p[1][13] , \p[1][12] , \p[1][11] , \p[0][28] , \p[0][27] ,
         \p[0][26] , \p[0][25] , \p[0][24] , \p[0][23] , \p[0][22] , \g[4][2] ,
         \g[3][2] , \g[2][6] , \g[2][5] , \g[1][13] , \g[1][12] , \g[1][11] ,
         \g[1][10] , \g[0][28] , \g[0][27] , \g[0][26] , \g[0][25] ,
         \g[0][24] , \g[0][23] , \g[0][22] , \g[0][21] ;

  PG_NETWORK_364 Block_PG_NET_21 ( .op1(A[20]), .op2(B[20]), .g(\g[0][21] ) );
  PG_NETWORK_363 Block_PG_NET_22 ( .op1(A[21]), .op2(B[21]), .g(\g[0][22] ), 
        .p(\p[0][22] ) );
  PG_NETWORK_362 Block_PG_NET_23 ( .op1(A[22]), .op2(B[22]), .g(\g[0][23] ), 
        .p(\p[0][23] ) );
  PG_NETWORK_361 Block_PG_NET_24 ( .op1(A[23]), .op2(B[23]), .g(\g[0][24] ), 
        .p(\p[0][24] ) );
  PG_NETWORK_360 Block_PG_NET_25 ( .op1(A[24]), .op2(B[24]), .g(\g[0][25] ), 
        .p(\p[0][25] ) );
  PG_NETWORK_359 Block_PG_NET_26 ( .op1(A[25]), .op2(B[25]), .g(\g[0][26] ), 
        .p(\p[0][26] ) );
  PG_NETWORK_358 Block_PG_NET_27 ( .op1(A[26]), .op2(B[26]), .g(\g[0][27] ), 
        .p(\p[0][27] ) );
  PG_NETWORK_357 Block_PG_NET_28 ( .op1(A[27]), .op2(B[27]), .g(\g[0][28] ), 
        .p(\p[0][28] ) );
  PG_BLOCK_369 Block_Stage_ONE_10 ( .P_ik(\p[0][22] ), .G_ik(\g[0][22] ), 
        .P_k1j(1'b0), .G_k1j(\g[0][21] ), .G_ij(\g[1][10] ) );
  PG_BLOCK_368 Block_Stage_ONE_11 ( .P_ik(\p[0][24] ), .G_ik(\g[0][24] ), 
        .P_k1j(\p[0][23] ), .G_k1j(\g[0][23] ), .P_ij(\p[1][11] ), .G_ij(
        \g[1][11] ) );
  PG_BLOCK_367 Block_Stage_ONE_12 ( .P_ik(\p[0][26] ), .G_ik(\g[0][26] ), 
        .P_k1j(\p[0][25] ), .G_k1j(\g[0][25] ), .P_ij(\p[1][12] ), .G_ij(
        \g[1][12] ) );
  PG_BLOCK_366 Block_Stage_ONE_13 ( .P_ik(\p[0][28] ), .G_ik(\g[0][28] ), 
        .P_k1j(\p[0][27] ), .G_k1j(\g[0][27] ), .P_ij(\p[1][13] ), .G_ij(
        \g[1][13] ) );
  PG_BLOCK_343 Block_Stage_TWO_5 ( .P_ik(\p[1][11] ), .G_ik(\g[1][11] ), 
        .P_k1j(1'b0), .G_k1j(\g[1][10] ), .G_ij_BAR(\g[2][5] ) );
  PG_BLOCK_342 Block_Stage_TWO_6 ( .P_ik(\p[1][13] ), .G_ik(\g[1][13] ), 
        .P_k1j(\p[1][12] ), .G_k1j(\g[1][12] ), .P_ij(\p[2][6] ), .G_ij(
        \g[2][6] ) );
  PG_BLOCK_331 Block_Stage_THREE_2 ( .P_ik(1'b0), .P_k1j(1'b0), .G_k1j(1'b0), 
        .G_ij_BAR(\g[3][2] ), .G_ik_BAR(\g[2][5] ) );
  PG_BLOCK_325 Block_stage_FOUR_2_0 ( .P_ik(\p[2][6] ), .G_ik(\g[2][6] ), 
        .P_k1j(1'b0), .G_ij_BAR(\g[4][2] ), .G_k1j_BAR(\g[3][2] ) );
  G_BLOCK_96 Block_stage_FIVE_5 ( .P_ik(1'b0), .G_k1j(1'b0), .G_ij(Cout[6]), 
        .G_ik_BAR(\g[3][2] ) );
  G_BLOCK_95 Block_stage_FIVE_6 ( .P_ik(1'b0), .G_k1j(1'b0), .G_ij(Cout[7]), 
        .G_ik_BAR(\g[4][2] ) );
endmodule


module FA_768 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_767 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_766 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_765 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_192 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_768 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_767 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_766 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_765 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_96 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_96 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_192 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0)
         );
  MUX_2to1_N4_96 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_760 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_759 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_758 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_757 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_190 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_760 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_759 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_758 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_757 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_95 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_95 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_190 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0)
         );
  MUX_2to1_N4_95 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_752 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_751 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_750 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_749 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_188 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_752 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_751 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_750 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_749 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_94 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_94 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_188 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0)
         );
  MUX_2to1_N4_94 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_744 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_743 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_742 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_741 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_186 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_744 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_743 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_742 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_741 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_93 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_93 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_186 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0)
         );
  MUX_2to1_N4_93 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_736 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_735 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_734 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_733 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_184 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_736 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_735 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_734 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_733 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_92 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_92 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_184 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0)
         );
  MUX_2to1_N4_92 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_728 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_727 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_726 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_725 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_182 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_728 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_727 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_726 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_725 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_91 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_91 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_182 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  MUX_2to1_N4_91 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_720 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_719 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_718 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_717 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_180 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_720 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_719 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_718 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_717 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_716 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_715 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_714 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_713 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_179 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_716 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_715 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_714 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_713 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_90 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U3 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U4 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
endmodule


module carry_select_block_N4_90 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_180 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_179 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_90 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_712 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_711 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_710 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_709 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_178 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_712 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_711 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_710 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_709 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_708 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_707 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_706 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_705 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_177 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_708 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_707 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_706 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_705 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_89 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U3 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U4 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
endmodule


module carry_select_block_N4_89 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_178 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_177 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_89 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module SUMGENERATOR_Nblocks16_bits_per_block4_6 ( A, B, CARRY_SELECT, SUM );
  input [63:0] A;
  input [63:0] B;
  input [15:0] CARRY_SELECT;
  output [63:0] SUM;


  carry_select_block_N4_96 block_n_1 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B[3:0]), .S(SUM[3:0]), .Ci(1'b0) );
  carry_select_block_N4_95 block_n_2 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B[7:4]), .S(SUM[7:4]), .Ci(1'b0) );
  carry_select_block_N4_94 block_n_3 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(
        B[11:8]), .S(SUM[11:8]), .Ci(1'b0) );
  carry_select_block_N4_93 block_n_4 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(
        B[15:12]), .S(SUM[15:12]), .Ci(1'b0) );
  carry_select_block_N4_92 block_n_5 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(
        B[19:16]), .S(SUM[19:16]), .Ci(1'b0) );
  carry_select_block_N4_91 block_n_6 ( .A(A[23:20]), .B(B[23:20]), .S(
        SUM[23:20]), .Ci(1'b0) );
  carry_select_block_N4_90 block_n_7 ( .A(A[27:24]), .B(B[27:24]), .S(
        SUM[27:24]), .Ci(CARRY_SELECT[6]) );
  carry_select_block_N4_89 block_n_8 ( .A(A[31:28]), .B(B[31:28]), .S(
        SUM[31:28]), .Ci(CARRY_SELECT[7]) );
endmodule


module ADDER_P4_N_BIT64_6 ( A, B, add_sub, Cout, SUM );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input add_sub;
  output Cout;

  wire   [63:0] B_xor;
  wire   [15:0] tmp_co;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46;
  assign B_xor[31] = B[31];
  assign B_xor[30] = B[30];
  assign B_xor[29] = B[29];
  assign B_xor[28] = B[28];
  assign B_xor[27] = B[27];
  assign B_xor[26] = B[26];
  assign B_xor[25] = B[25];
  assign B_xor[24] = B[24];
  assign B_xor[23] = B[23];
  assign B_xor[22] = B[22];
  assign B_xor[21] = B[21];
  assign B_xor[20] = B[20];
  assign B_xor[19] = B[19];
  assign B_xor[18] = B[18];
  assign B_xor[17] = B[17];
  assign B_xor[16] = B[16];
  assign B_xor[15] = B[15];
  assign B_xor[14] = B[14];
  assign B_xor[13] = B[13];
  assign B_xor[12] = B[12];
  assign B_xor[11] = B[11];
  assign B_xor[10] = B[10];
  assign B_xor[9] = B[9];
  assign B_xor[8] = B[8];
  assign B_xor[7] = B[7];
  assign B_xor[6] = B[6];
  assign B_xor[5] = B[5];
  assign B_xor[4] = B[4];
  assign B_xor[3] = B[3];
  assign B_xor[2] = B[2];
  assign B_xor[1] = B[1];
  assign B_xor[0] = B[0];

  CARRY_GENERATOR_Nbit64_6 CLA_SPARSE_TREE ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, A[27:20], 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B_xor[27:20], 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Cin(1'b0), .Cout({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, tmp_co[7:6], SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14}) );
  SUMGENERATOR_Nblocks16_bits_per_block4_6 CSA ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, A[31:20], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        B_xor[31:0]}), .CARRY_SELECT({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, tmp_co[7:6], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .SUM({
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, SYNOPSYS_UNCONNECTED__22, 
        SYNOPSYS_UNCONNECTED__23, SYNOPSYS_UNCONNECTED__24, 
        SYNOPSYS_UNCONNECTED__25, SYNOPSYS_UNCONNECTED__26, 
        SYNOPSYS_UNCONNECTED__27, SYNOPSYS_UNCONNECTED__28, 
        SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, 
        SYNOPSYS_UNCONNECTED__31, SYNOPSYS_UNCONNECTED__32, 
        SYNOPSYS_UNCONNECTED__33, SYNOPSYS_UNCONNECTED__34, 
        SYNOPSYS_UNCONNECTED__35, SYNOPSYS_UNCONNECTED__36, 
        SYNOPSYS_UNCONNECTED__37, SYNOPSYS_UNCONNECTED__38, 
        SYNOPSYS_UNCONNECTED__39, SYNOPSYS_UNCONNECTED__40, 
        SYNOPSYS_UNCONNECTED__41, SYNOPSYS_UNCONNECTED__42, 
        SYNOPSYS_UNCONNECTED__43, SYNOPSYS_UNCONNECTED__44, 
        SYNOPSYS_UNCONNECTED__45, SYNOPSYS_UNCONNECTED__46, SUM[31:0]}) );
endmodule


module PG_NETWORK_298 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_297 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_296 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_295 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_294 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_293 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_BLOCK_305 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij_BAR );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij_BAR;


  AOI21_X1 U1 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(G_ij_BAR) );
endmodule


module PG_BLOCK_304 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_303 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_280 ( P_ik, P_k1j, G_k1j, P_ij, G_ij_BAR, G_ik_BAR );
  input P_ik, P_k1j, G_k1j, G_ik_BAR;
  output P_ij, G_ij_BAR;
  wire   G_ik;
  assign G_ij_BAR = G_ik;
  assign G_ik = G_ik_BAR;

endmodule


module PG_BLOCK_279 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_268 ( P_ik, P_k1j, G_k1j, P_ij, G_ij_BAR, G_ik_BAR );
  input P_ik, P_k1j, G_k1j, G_ik_BAR;
  output P_ij, G_ij_BAR;
  wire   G_ik;
  assign G_ij_BAR = G_ik;
  assign G_ik = G_ik_BAR;

endmodule


module PG_BLOCK_262 ( P_ik, G_ik, P_k1j, P_ij, G_ij_BAR, G_k1j_BAR );
  input P_ik, G_ik, P_k1j, G_k1j_BAR;
  output P_ij, G_ij_BAR;
  wire   G_k1j, n1;
  assign G_k1j = G_k1j_BAR;

  INV_X1 U1 ( .A(G_k1j), .ZN(n1) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(n1), .A(G_ik), .ZN(G_ij_BAR) );
endmodule


module G_BLOCK_79 ( P_ik, G_k1j, G_ij, G_ik_BAR );
  input P_ik, G_k1j, G_ik_BAR;
  output G_ij;
  wire   G_ik;
  assign G_ik = G_ik_BAR;

  INV_X1 U1 ( .A(G_ik), .ZN(G_ij) );
endmodule


module G_BLOCK_78 ( P_ik, G_k1j, G_ij, G_ik_BAR );
  input P_ik, G_k1j, G_ik_BAR;
  output G_ij;
  wire   G_ik;
  assign G_ik = G_ik_BAR;

  INV_X1 U1 ( .A(G_ik), .ZN(G_ij) );
endmodule


module CARRY_GENERATOR_Nbit64_5 ( A, B, Cin, Cout );
  input [63:0] A;
  input [63:0] B;
  output [16:0] Cout;
  input Cin;
  wire   \p[2][6] , \p[1][13] , \p[1][12] , \p[0][28] , \p[0][27] , \p[0][26] ,
         \p[0][25] , \p[0][24] , \g[4][2] , \g[3][2] , \g[2][6] , \g[2][5] ,
         \g[1][13] , \g[1][12] , \g[1][11] , \g[0][28] , \g[0][27] ,
         \g[0][26] , \g[0][25] , \g[0][24] , \g[0][23] ;

  PG_NETWORK_298 Block_PG_NET_23 ( .op1(A[22]), .op2(B[22]), .g(\g[0][23] ) );
  PG_NETWORK_297 Block_PG_NET_24 ( .op1(A[23]), .op2(B[23]), .g(\g[0][24] ), 
        .p(\p[0][24] ) );
  PG_NETWORK_296 Block_PG_NET_25 ( .op1(A[24]), .op2(B[24]), .g(\g[0][25] ), 
        .p(\p[0][25] ) );
  PG_NETWORK_295 Block_PG_NET_26 ( .op1(A[25]), .op2(B[25]), .g(\g[0][26] ), 
        .p(\p[0][26] ) );
  PG_NETWORK_294 Block_PG_NET_27 ( .op1(A[26]), .op2(B[26]), .g(\g[0][27] ), 
        .p(\p[0][27] ) );
  PG_NETWORK_293 Block_PG_NET_28 ( .op1(A[27]), .op2(B[27]), .g(\g[0][28] ), 
        .p(\p[0][28] ) );
  PG_BLOCK_305 Block_Stage_ONE_11 ( .P_ik(\p[0][24] ), .G_ik(\g[0][24] ), 
        .P_k1j(1'b0), .G_k1j(\g[0][23] ), .G_ij_BAR(\g[1][11] ) );
  PG_BLOCK_304 Block_Stage_ONE_12 ( .P_ik(\p[0][26] ), .G_ik(\g[0][26] ), 
        .P_k1j(\p[0][25] ), .G_k1j(\g[0][25] ), .P_ij(\p[1][12] ), .G_ij(
        \g[1][12] ) );
  PG_BLOCK_303 Block_Stage_ONE_13 ( .P_ik(\p[0][28] ), .G_ik(\g[0][28] ), 
        .P_k1j(\p[0][27] ), .G_k1j(\g[0][27] ), .P_ij(\p[1][13] ), .G_ij(
        \g[1][13] ) );
  PG_BLOCK_280 Block_Stage_TWO_5 ( .P_ik(1'b0), .P_k1j(1'b0), .G_k1j(1'b0), 
        .G_ij_BAR(\g[2][5] ), .G_ik_BAR(\g[1][11] ) );
  PG_BLOCK_279 Block_Stage_TWO_6 ( .P_ik(\p[1][13] ), .G_ik(\g[1][13] ), 
        .P_k1j(\p[1][12] ), .G_k1j(\g[1][12] ), .P_ij(\p[2][6] ), .G_ij(
        \g[2][6] ) );
  PG_BLOCK_268 Block_Stage_THREE_2 ( .P_ik(1'b0), .P_k1j(1'b0), .G_k1j(1'b0), 
        .G_ij_BAR(\g[3][2] ), .G_ik_BAR(\g[2][5] ) );
  PG_BLOCK_262 Block_stage_FOUR_2_0 ( .P_ik(\p[2][6] ), .G_ik(\g[2][6] ), 
        .P_k1j(1'b0), .G_ij_BAR(\g[4][2] ), .G_k1j_BAR(\g[3][2] ) );
  G_BLOCK_79 Block_stage_FIVE_5 ( .P_ik(1'b0), .G_k1j(1'b0), .G_ij(Cout[6]), 
        .G_ik_BAR(\g[3][2] ) );
  G_BLOCK_78 Block_stage_FIVE_6 ( .P_ik(1'b0), .G_k1j(1'b0), .G_ij(Cout[7]), 
        .G_ik_BAR(\g[4][2] ) );
endmodule


module FA_640 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_639 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_638 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_637 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_160 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_640 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_639 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_638 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_637 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_80 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_80 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_160 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0)
         );
  MUX_2to1_N4_80 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_632 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_631 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_630 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_629 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_158 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_632 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_631 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_630 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_629 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_79 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_79 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_158 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0)
         );
  MUX_2to1_N4_79 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_624 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_623 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_622 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_621 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_156 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_624 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_623 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_622 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_621 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_78 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_78 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_156 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0)
         );
  MUX_2to1_N4_78 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_616 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_615 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_614 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_613 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_154 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_616 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_615 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_614 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_613 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_77 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_77 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_154 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0)
         );
  MUX_2to1_N4_77 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_608 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_607 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_606 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_605 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_152 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_608 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_607 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_606 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_605 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_76 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_76 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_152 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0)
         );
  MUX_2to1_N4_76 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_600 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_599 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_598 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_597 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_150 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \CTMP[3] ;

  FA_600 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_599 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_598 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(1'b0), .S(S[2]), .Co(\CTMP[3] )
         );
  FA_597 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(\CTMP[3] ), .S(S[3]) );
endmodule


module MUX_2to1_N4_75 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_75 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_150 RCA_0 ( .A({A[3:2], 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0) );
  MUX_2to1_N4_75 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_592 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_591 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_590 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_589 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_148 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_592 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_591 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_590 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_589 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_588 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_587 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_586 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_585 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_147 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_588 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_587 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_586 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_585 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_74 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U3 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U4 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
endmodule


module carry_select_block_N4_74 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_148 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_147 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_74 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module FA_584 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_583 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_582 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_581 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_146 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_584 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_583 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_582 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_581 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_580 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_579 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_578 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_577 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_145 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_580 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_579 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_578 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_577 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_73 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U3 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U4 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
endmodule


module carry_select_block_N4_73 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_146 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_145 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_73 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module SUMGENERATOR_Nblocks16_bits_per_block4_5 ( A, B, CARRY_SELECT, SUM );
  input [63:0] A;
  input [63:0] B;
  input [15:0] CARRY_SELECT;
  output [63:0] SUM;


  carry_select_block_N4_80 block_n_1 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B[3:0]), .S(SUM[3:0]), .Ci(1'b0) );
  carry_select_block_N4_79 block_n_2 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B[7:4]), .S(SUM[7:4]), .Ci(1'b0) );
  carry_select_block_N4_78 block_n_3 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(
        B[11:8]), .S(SUM[11:8]), .Ci(1'b0) );
  carry_select_block_N4_77 block_n_4 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(
        B[15:12]), .S(SUM[15:12]), .Ci(1'b0) );
  carry_select_block_N4_76 block_n_5 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(
        B[19:16]), .S(SUM[19:16]), .Ci(1'b0) );
  carry_select_block_N4_75 block_n_6 ( .A({A[23:22], 1'b0, 1'b0}), .B(B[23:20]), .S(SUM[23:20]), .Ci(1'b0) );
  carry_select_block_N4_74 block_n_7 ( .A(A[27:24]), .B(B[27:24]), .S(
        SUM[27:24]), .Ci(CARRY_SELECT[6]) );
  carry_select_block_N4_73 block_n_8 ( .A(A[31:28]), .B(B[31:28]), .S(
        SUM[31:28]), .Ci(CARRY_SELECT[7]) );
endmodule


module ADDER_P4_N_BIT64_5 ( A, B, add_sub, Cout, SUM );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input add_sub;
  output Cout;

  wire   [63:0] B_xor;
  wire   [15:0] tmp_co;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46;
  assign B_xor[31] = B[31];
  assign B_xor[30] = B[30];
  assign B_xor[29] = B[29];
  assign B_xor[28] = B[28];
  assign B_xor[27] = B[27];
  assign B_xor[26] = B[26];
  assign B_xor[25] = B[25];
  assign B_xor[24] = B[24];
  assign B_xor[23] = B[23];
  assign B_xor[22] = B[22];
  assign B_xor[21] = B[21];
  assign B_xor[20] = B[20];
  assign B_xor[19] = B[19];
  assign B_xor[18] = B[18];
  assign B_xor[17] = B[17];
  assign B_xor[16] = B[16];
  assign B_xor[15] = B[15];
  assign B_xor[14] = B[14];
  assign B_xor[13] = B[13];
  assign B_xor[12] = B[12];
  assign B_xor[11] = B[11];
  assign B_xor[10] = B[10];
  assign B_xor[9] = B[9];
  assign B_xor[8] = B[8];
  assign B_xor[7] = B[7];
  assign B_xor[6] = B[6];
  assign B_xor[5] = B[5];
  assign B_xor[4] = B[4];
  assign B_xor[3] = B[3];
  assign B_xor[2] = B[2];
  assign B_xor[1] = B[1];
  assign B_xor[0] = B[0];

  CARRY_GENERATOR_Nbit64_5 CLA_SPARSE_TREE ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, A[27:22], 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B_xor[27:22], 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Cin(1'b0), 
        .Cout({SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, tmp_co[7:6], SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14}) );
  SUMGENERATOR_Nblocks16_bits_per_block4_5 CSA ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, A[31:22], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, B_xor[31:0]}), .CARRY_SELECT({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, tmp_co[7:6], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .SUM({
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, SYNOPSYS_UNCONNECTED__22, 
        SYNOPSYS_UNCONNECTED__23, SYNOPSYS_UNCONNECTED__24, 
        SYNOPSYS_UNCONNECTED__25, SYNOPSYS_UNCONNECTED__26, 
        SYNOPSYS_UNCONNECTED__27, SYNOPSYS_UNCONNECTED__28, 
        SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, 
        SYNOPSYS_UNCONNECTED__31, SYNOPSYS_UNCONNECTED__32, 
        SYNOPSYS_UNCONNECTED__33, SYNOPSYS_UNCONNECTED__34, 
        SYNOPSYS_UNCONNECTED__35, SYNOPSYS_UNCONNECTED__36, 
        SYNOPSYS_UNCONNECTED__37, SYNOPSYS_UNCONNECTED__38, 
        SYNOPSYS_UNCONNECTED__39, SYNOPSYS_UNCONNECTED__40, 
        SYNOPSYS_UNCONNECTED__41, SYNOPSYS_UNCONNECTED__42, 
        SYNOPSYS_UNCONNECTED__43, SYNOPSYS_UNCONNECTED__44, 
        SYNOPSYS_UNCONNECTED__45, SYNOPSYS_UNCONNECTED__46, SUM[31:0]}) );
endmodule


module PG_NETWORK_232 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_231 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_230 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_NETWORK_229 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
  XOR2_X1 U2 ( .A(op2), .B(op1), .Z(p) );
endmodule


module PG_BLOCK_241 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AOI21_X1 U1 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_240 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij;
  wire   n1;

  AND2_X1 U1 ( .A1(P_ik), .A2(P_k1j), .ZN(P_ij) );
  AOI21_X1 U2 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(n1) );
  INV_X1 U3 ( .A(n1), .ZN(G_ij) );
endmodule


module PG_BLOCK_216 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij_BAR );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij_BAR;


  AOI21_X1 U1 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(G_ij_BAR) );
endmodule


module PG_BLOCK_199 ( P_ik, P_k1j, G_k1j, P_ij, G_ij_BAR, G_ik_BAR );
  input P_ik, P_k1j, G_k1j, G_ik_BAR;
  output P_ij, G_ij_BAR;
  wire   G_ik;
  assign G_ij_BAR = G_ik;
  assign G_ik = G_ik_BAR;

endmodule


module G_BLOCK_61 ( P_ik, G_k1j, G_ij, G_ik_BAR );
  input P_ik, G_k1j, G_ik_BAR;
  output G_ij;
  wire   G_ik;
  assign G_ik = G_ik_BAR;

  INV_X1 U1 ( .A(G_ik), .ZN(G_ij) );
endmodule


module CARRY_GENERATOR_Nbit64_4 ( A, B, Cin, Cout );
  input [63:0] A;
  input [63:0] B;
  output [16:0] Cout;
  input Cin;
  wire   \p[1][13] , \p[0][28] , \p[0][27] , \p[0][26] , \g[4][2] , \g[2][6] ,
         \g[1][13] , \g[1][12] , \g[0][28] , \g[0][27] , \g[0][26] ,
         \g[0][25] ;

  PG_NETWORK_232 Block_PG_NET_25 ( .op1(A[24]), .op2(B[24]), .g(\g[0][25] ) );
  PG_NETWORK_231 Block_PG_NET_26 ( .op1(A[25]), .op2(B[25]), .g(\g[0][26] ), 
        .p(\p[0][26] ) );
  PG_NETWORK_230 Block_PG_NET_27 ( .op1(A[26]), .op2(B[26]), .g(\g[0][27] ), 
        .p(\p[0][27] ) );
  PG_NETWORK_229 Block_PG_NET_28 ( .op1(A[27]), .op2(B[27]), .g(\g[0][28] ), 
        .p(\p[0][28] ) );
  PG_BLOCK_241 Block_Stage_ONE_12 ( .P_ik(\p[0][26] ), .G_ik(\g[0][26] ), 
        .P_k1j(1'b0), .G_k1j(\g[0][25] ), .G_ij(\g[1][12] ) );
  PG_BLOCK_240 Block_Stage_ONE_13 ( .P_ik(\p[0][28] ), .G_ik(\g[0][28] ), 
        .P_k1j(\p[0][27] ), .G_k1j(\g[0][27] ), .P_ij(\p[1][13] ), .G_ij(
        \g[1][13] ) );
  PG_BLOCK_216 Block_Stage_TWO_6 ( .P_ik(\p[1][13] ), .G_ik(\g[1][13] ), 
        .P_k1j(1'b0), .G_k1j(\g[1][12] ), .G_ij_BAR(\g[2][6] ) );
  PG_BLOCK_199 Block_stage_FOUR_2_0 ( .P_ik(1'b0), .P_k1j(1'b0), .G_k1j(1'b0), 
        .G_ij_BAR(\g[4][2] ), .G_ik_BAR(\g[2][6] ) );
  G_BLOCK_61 Block_stage_FIVE_6 ( .P_ik(1'b0), .G_k1j(1'b0), .G_ij(Cout[7]), 
        .G_ik_BAR(\g[4][2] ) );
endmodule


module FA_512 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_511 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_510 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_509 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_128 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_512 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_511 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_510 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_509 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_64 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_64 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_128 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0)
         );
  MUX_2to1_N4_64 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_504 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_503 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_502 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_501 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_126 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_504 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_503 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_502 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_501 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_63 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_63 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_126 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0)
         );
  MUX_2to1_N4_63 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_496 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_495 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_494 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_493 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_124 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_496 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_495 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_494 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_493 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_62 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_62 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_124 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0)
         );
  MUX_2to1_N4_62 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_488 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_487 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_486 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_485 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_122 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_488 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_487 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_486 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_485 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_61 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_61 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_122 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0)
         );
  MUX_2to1_N4_61 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_480 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_479 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_478 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_477 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_120 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_480 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_479 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_478 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_477 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_60 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_60 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_120 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0)
         );
  MUX_2to1_N4_60 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_472 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_471 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_470 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_469 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_118 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_472 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_471 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_470 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_469 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_59 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_59 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_118 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0)
         );
  MUX_2to1_N4_59 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_464 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_463 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_462 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_461 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_116 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_464 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_463 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_462 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_461 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_58 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_58 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_116 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  MUX_2to1_N4_58 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_456 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_455 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_454 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_453 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_114 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_456 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_455 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_454 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_453 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_452 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_451 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_450 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_449 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_113 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_452 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_451 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_450 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_449 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_57 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;


  MUX2_X1 U1 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U3 ( .A(IN0[2]), .B(IN1[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U4 ( .A(IN0[3]), .B(IN1[3]), .S(SEL), .Z(Y[3]) );
endmodule


module carry_select_block_N4_57 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_114 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_113 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_57 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module SUMGENERATOR_Nblocks16_bits_per_block4_4 ( A, B, CARRY_SELECT, SUM );
  input [63:0] A;
  input [63:0] B;
  input [15:0] CARRY_SELECT;
  output [63:0] SUM;


  carry_select_block_N4_64 block_n_1 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B[3:0]), .S(SUM[3:0]), .Ci(1'b0) );
  carry_select_block_N4_63 block_n_2 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B[7:4]), .S(SUM[7:4]), .Ci(1'b0) );
  carry_select_block_N4_62 block_n_3 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(
        B[11:8]), .S(SUM[11:8]), .Ci(1'b0) );
  carry_select_block_N4_61 block_n_4 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(
        B[15:12]), .S(SUM[15:12]), .Ci(1'b0) );
  carry_select_block_N4_60 block_n_5 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(
        B[19:16]), .S(SUM[19:16]), .Ci(1'b0) );
  carry_select_block_N4_59 block_n_6 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(
        B[23:20]), .S(SUM[23:20]), .Ci(1'b0) );
  carry_select_block_N4_58 block_n_7 ( .A(A[27:24]), .B(B[27:24]), .S(
        SUM[27:24]), .Ci(1'b0) );
  carry_select_block_N4_57 block_n_8 ( .A(A[31:28]), .B(B[31:28]), .S(
        SUM[31:28]), .Ci(CARRY_SELECT[7]) );
endmodule


module ADDER_P4_N_BIT64_4 ( A, B, add_sub, Cout, SUM );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input add_sub;
  output Cout;
  wire   \tmp_co[7] ;
  wire   [63:0] B_xor;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47;
  assign B_xor[31] = B[31];
  assign B_xor[30] = B[30];
  assign B_xor[29] = B[29];
  assign B_xor[28] = B[28];
  assign B_xor[27] = B[27];
  assign B_xor[26] = B[26];
  assign B_xor[25] = B[25];
  assign B_xor[24] = B[24];
  assign B_xor[23] = B[23];
  assign B_xor[22] = B[22];
  assign B_xor[21] = B[21];
  assign B_xor[20] = B[20];
  assign B_xor[19] = B[19];
  assign B_xor[18] = B[18];
  assign B_xor[17] = B[17];
  assign B_xor[16] = B[16];
  assign B_xor[15] = B[15];
  assign B_xor[14] = B[14];
  assign B_xor[13] = B[13];
  assign B_xor[12] = B[12];
  assign B_xor[11] = B[11];
  assign B_xor[10] = B[10];
  assign B_xor[9] = B[9];
  assign B_xor[8] = B[8];
  assign B_xor[7] = B[7];
  assign B_xor[6] = B[6];
  assign B_xor[5] = B[5];
  assign B_xor[4] = B[4];
  assign B_xor[3] = B[3];
  assign B_xor[2] = B[2];
  assign B_xor[1] = B[1];
  assign B_xor[0] = B[0];

  CARRY_GENERATOR_Nbit64_4 CLA_SPARSE_TREE ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, A[27:24], 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        B_xor[27:24], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .Cin(1'b0), .Cout({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, \tmp_co[7] , 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15}) );
  SUMGENERATOR_Nblocks16_bits_per_block4_4 CSA ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, A[31:24], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, B_xor[31:0]}), .CARRY_SELECT({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, \tmp_co[7] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .SUM({SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, SUM[31:0]}) );
endmodule


module PG_NETWORK_166 ( op1, op2, g, p );
  input op1, op2;
  output g, p;


  AND2_X1 U1 ( .A1(op2), .A2(op1), .ZN(g) );
endmodule


module PG_NETWORK_165 ( op1, op2, g, p );
  input op1, op2;
  output g, p;
  wire   n1;

  XNOR2_X1 U1 ( .A(op1), .B(n1), .ZN(p) );
  INV_X1 U2 ( .A(op2), .ZN(n1) );
  AND2_X1 U3 ( .A1(op1), .A2(op2), .ZN(g) );
endmodule


module PG_BLOCK_177 ( P_ik, G_ik, P_k1j, G_k1j, P_ij, G_ij_BAR );
  input P_ik, G_ik, P_k1j, G_k1j;
  output P_ij, G_ij_BAR;


  AOI21_X1 U1 ( .B1(G_k1j), .B2(P_ik), .A(G_ik), .ZN(G_ij_BAR) );
endmodule


module PG_BLOCK_153 ( P_ik, P_k1j, G_k1j, P_ij, G_ij_BAR, G_ik_BAR );
  input P_ik, P_k1j, G_k1j, G_ik_BAR;
  output P_ij, G_ij_BAR;
  wire   G_ik;
  assign G_ij_BAR = G_ik;
  assign G_ik = G_ik_BAR;

endmodule


module PG_BLOCK_136 ( P_ik, P_k1j, G_k1j, P_ij, G_ij_BAR, G_ik_BAR );
  input P_ik, P_k1j, G_k1j, G_ik_BAR;
  output P_ij, G_ij_BAR;
  wire   G_ik;
  assign G_ij_BAR = G_ik;
  assign G_ik = G_ik_BAR;

endmodule


module G_BLOCK_44 ( P_ik, G_k1j, G_ij, G_ik_BAR );
  input P_ik, G_k1j, G_ik_BAR;
  output G_ij;
  wire   G_ik;
  assign G_ik = G_ik_BAR;

  INV_X1 U1 ( .A(G_ik), .ZN(G_ij) );
endmodule


module CARRY_GENERATOR_Nbit64_3 ( A, B, Cin, Cout );
  input [63:0] A;
  input [63:0] B;
  output [16:0] Cout;
  input Cin;
  wire   \p[0][28] , \g[4][2] , \g[2][6] , \g[1][13] , \g[0][28] , \g[0][27] ;

  PG_NETWORK_166 Block_PG_NET_27 ( .op1(A[26]), .op2(B[26]), .g(\g[0][27] ) );
  PG_NETWORK_165 Block_PG_NET_28 ( .op1(A[27]), .op2(B[27]), .g(\g[0][28] ), 
        .p(\p[0][28] ) );
  PG_BLOCK_177 Block_Stage_ONE_13 ( .P_ik(\p[0][28] ), .G_ik(\g[0][28] ), 
        .P_k1j(1'b0), .G_k1j(\g[0][27] ), .G_ij_BAR(\g[1][13] ) );
  PG_BLOCK_153 Block_Stage_TWO_6 ( .P_ik(1'b0), .P_k1j(1'b0), .G_k1j(1'b0), 
        .G_ij_BAR(\g[2][6] ), .G_ik_BAR(\g[1][13] ) );
  PG_BLOCK_136 Block_stage_FOUR_2_0 ( .P_ik(1'b0), .P_k1j(1'b0), .G_k1j(1'b0), 
        .G_ij_BAR(\g[4][2] ), .G_ik_BAR(\g[2][6] ) );
  G_BLOCK_44 Block_stage_FIVE_6 ( .P_ik(1'b0), .G_k1j(1'b0), .G_ij(Cout[7]), 
        .G_ik_BAR(\g[4][2] ) );
endmodule


module FA_384 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_383 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_382 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_381 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_96 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_384 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_383 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_382 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_381 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_48 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_48 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_96 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0) );
  MUX_2to1_N4_48 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_376 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_375 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_374 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_373 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_94 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_376 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_375 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_374 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_373 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_47 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_47 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_94 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0) );
  MUX_2to1_N4_47 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_368 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_367 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_366 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_365 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_92 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_368 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_367 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_366 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_365 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_46 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_46 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_92 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0) );
  MUX_2to1_N4_46 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_360 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_359 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_358 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_357 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_90 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_360 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_359 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_358 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_357 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_45 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_45 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_90 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0) );
  MUX_2to1_N4_45 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_352 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_351 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_350 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_349 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_88 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_352 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_351 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_350 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_349 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_44 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_44 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_88 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0) );
  MUX_2to1_N4_44 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_344 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_343 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_342 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_341 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_86 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_344 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_343 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_342 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_341 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_43 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_43 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_86 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0) );
  MUX_2to1_N4_43 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_336 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_335 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_334 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_333 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_84 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \CTMP[3] ;

  FA_336 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_335 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_334 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(1'b0), .S(S[2]), .Co(\CTMP[3] )
         );
  FA_333 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(\CTMP[3] ), .S(S[3]) );
endmodule


module MUX_2to1_N4_42 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_42 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_84 RCA_0 ( .A({A[3:2], 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0) );
  MUX_2to1_N4_42 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_328 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_327 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_326 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_325 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_82 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_328 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_327 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_326 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_325 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module FA_324 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  OR2_X1 U1 ( .A1(A), .A2(B), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(S) );
endmodule


module FA_323 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4;

  XNOR2_X1 U1 ( .A(Ci), .B(n4), .ZN(S) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n2), .A2(n1), .ZN(Co) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n1) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n3), .ZN(n2) );
  OR2_X1 U6 ( .A1(A), .A2(B), .ZN(n3) );
endmodule


module FA_322 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_321 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_81 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_324 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b1), .S(S[0]), .Co(CTMP[1])
         );
  FA_323 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_322 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_321 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_41 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;
  wire   n1, n2, n3, n4;

  NAND2_X1 U1 ( .A1(n1), .A2(n3), .ZN(Y[3]) );
  NAND2_X1 U2 ( .A1(IN0[3]), .A2(n2), .ZN(n1) );
  INV_X1 U3 ( .A(n4), .ZN(n2) );
  NAND2_X1 U4 ( .A1(IN1[3]), .A2(n4), .ZN(n3) );
  BUF_X1 U5 ( .A(SEL), .Z(n4) );
  MUX2_X1 U6 ( .A(IN0[0]), .B(IN1[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U7 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U8 ( .A(IN0[2]), .B(IN1[2]), .S(n4), .Z(Y[2]) );
endmodule


module carry_select_block_N4_41 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;
  wire   [3:0] S_1;

  RCA_N4_82 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  RCA_N4_81 RCA_1 ( .A(A), .B(B), .Ci(1'b1), .S(S_1) );
  MUX_2to1_N4_41 SUM_SELECT_MUX ( .IN0(S_0), .IN1(S_1), .SEL(Ci), .Y(S) );
endmodule


module SUMGENERATOR_Nblocks16_bits_per_block4_3 ( A, B, CARRY_SELECT, SUM );
  input [63:0] A;
  input [63:0] B;
  input [15:0] CARRY_SELECT;
  output [63:0] SUM;


  carry_select_block_N4_48 block_n_1 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B[3:0]), .S(SUM[3:0]), .Ci(1'b0) );
  carry_select_block_N4_47 block_n_2 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B[7:4]), .S(SUM[7:4]), .Ci(1'b0) );
  carry_select_block_N4_46 block_n_3 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(
        B[11:8]), .S(SUM[11:8]), .Ci(1'b0) );
  carry_select_block_N4_45 block_n_4 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(
        B[15:12]), .S(SUM[15:12]), .Ci(1'b0) );
  carry_select_block_N4_44 block_n_5 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(
        B[19:16]), .S(SUM[19:16]), .Ci(1'b0) );
  carry_select_block_N4_43 block_n_6 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(
        B[23:20]), .S(SUM[23:20]), .Ci(1'b0) );
  carry_select_block_N4_42 block_n_7 ( .A({A[27:26], 1'b0, 1'b0}), .B(B[27:24]), .S(SUM[27:24]), .Ci(1'b0) );
  carry_select_block_N4_41 block_n_8 ( .A(A[31:28]), .B(B[31:28]), .S(
        SUM[31:28]), .Ci(CARRY_SELECT[7]) );
endmodule


module ADDER_P4_N_BIT64_3 ( A, B, add_sub, Cout, SUM );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input add_sub;
  output Cout;
  wire   \tmp_co[7] , n1;
  wire   [63:0] B_xor;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47;
  assign B_xor[31] = B[31];
  assign B_xor[30] = B[30];
  assign B_xor[29] = B[29];
  assign B_xor[28] = B[28];
  assign B_xor[27] = B[27];
  assign B_xor[26] = B[26];
  assign B_xor[25] = B[25];
  assign B_xor[24] = B[24];
  assign B_xor[23] = B[23];
  assign B_xor[22] = B[22];
  assign B_xor[21] = B[21];
  assign B_xor[20] = B[20];
  assign B_xor[19] = B[19];
  assign B_xor[18] = B[18];
  assign B_xor[17] = B[17];
  assign B_xor[16] = B[16];
  assign B_xor[15] = B[15];
  assign B_xor[14] = B[14];
  assign B_xor[13] = B[13];
  assign B_xor[12] = B[12];
  assign B_xor[11] = B[11];
  assign B_xor[10] = B[10];
  assign B_xor[9] = B[9];
  assign B_xor[8] = B[8];
  assign B_xor[7] = B[7];
  assign B_xor[6] = B[6];
  assign B_xor[5] = B[5];
  assign B_xor[4] = B[4];
  assign B_xor[3] = B[3];
  assign B_xor[2] = B[2];
  assign B_xor[1] = B[1];
  assign B_xor[0] = B[0];

  CARRY_GENERATOR_Nbit64_3 CLA_SPARSE_TREE ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, A[27:26], 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, B_xor[27:26], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Cin(1'b0), .Cout({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, \tmp_co[7] , SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15}) );
  SUMGENERATOR_Nblocks16_bits_per_block4_3 CSA ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, A[31:28], n1, A[26], 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B_xor[31:0]}), 
        .CARRY_SELECT({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        \tmp_co[7] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .SUM({
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, SUM[31:0]}) );
  BUF_X1 U1 ( .A(A[27]), .Z(n1) );
endmodule


module FA_256 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_255 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_254 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_253 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_64 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_256 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_255 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_254 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_253 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_32 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_32 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_64 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0) );
  MUX_2to1_N4_32 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_248 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_247 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_246 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_245 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_62 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_248 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_247 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_246 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_245 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_31 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_31 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_62 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0) );
  MUX_2to1_N4_31 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_240 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_239 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_238 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_237 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_60 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_240 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_239 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_238 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_237 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_30 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_30 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_60 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0) );
  MUX_2to1_N4_30 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_232 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_231 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_230 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_229 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_58 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_232 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_231 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_230 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_229 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_29 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_29 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_58 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0) );
  MUX_2to1_N4_29 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_224 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_223 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_222 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_221 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_56 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_224 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_223 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_222 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_221 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_28 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_28 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_56 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0) );
  MUX_2to1_N4_28 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_216 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_215 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_214 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_213 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_54 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_216 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_215 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_214 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_213 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_27 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_27 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_54 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0) );
  MUX_2to1_N4_27 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_208 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_207 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_206 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_205 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_52 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_208 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_207 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_206 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_205 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_26 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_26 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_52 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0) );
  MUX_2to1_N4_26 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_200 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(Co) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_199 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  FA_X1 U1 ( .A(A), .B(B), .CI(Ci), .CO(Co), .S(S) );
endmodule


module FA_198 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1, n2, n3, n4;

  BUF_X1 U1 ( .A(Ci), .Z(n1) );
  NAND2_X1 U2 ( .A1(B), .A2(A), .ZN(n3) );
  NAND2_X1 U3 ( .A1(n3), .A2(n2), .ZN(Co) );
  OAI21_X1 U4 ( .B1(A), .B2(B), .A(Ci), .ZN(n2) );
  XNOR2_X1 U5 ( .A(n4), .B(n1), .ZN(S) );
  XNOR2_X1 U6 ( .A(B), .B(A), .ZN(n4) );
endmodule


module FA_197 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n1) );
  XNOR2_X1 U2 ( .A(Ci), .B(n1), .ZN(S) );
endmodule


module RCA_N4_50 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_200 FULLADDER_1 ( .A(A[0]), .B(B[0]), .Ci(1'b0), .S(S[0]), .Co(CTMP[1])
         );
  FA_199 FULLADDER_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_198 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_197 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]) );
endmodule


module MUX_2to1_N4_25 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_25 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_50 RCA_0 ( .A(A), .B(B), .Ci(1'b0), .S(S_0) );
  MUX_2to1_N4_25 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module SUMGENERATOR_Nblocks16_bits_per_block4_2 ( A, B, CARRY_SELECT, SUM );
  input [63:0] A;
  input [63:0] B;
  input [15:0] CARRY_SELECT;
  output [63:0] SUM;


  carry_select_block_N4_32 block_n_1 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B[3:0]), .S(SUM[3:0]), .Ci(1'b0) );
  carry_select_block_N4_31 block_n_2 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B[7:4]), .S(SUM[7:4]), .Ci(1'b0) );
  carry_select_block_N4_30 block_n_3 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(
        B[11:8]), .S(SUM[11:8]), .Ci(1'b0) );
  carry_select_block_N4_29 block_n_4 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(
        B[15:12]), .S(SUM[15:12]), .Ci(1'b0) );
  carry_select_block_N4_28 block_n_5 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(
        B[19:16]), .S(SUM[19:16]), .Ci(1'b0) );
  carry_select_block_N4_27 block_n_6 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(
        B[23:20]), .S(SUM[23:20]), .Ci(1'b0) );
  carry_select_block_N4_26 block_n_7 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(
        B[27:24]), .S(SUM[27:24]), .Ci(1'b0) );
  carry_select_block_N4_25 block_n_8 ( .A(A[31:28]), .B(B[31:28]), .S(
        SUM[31:28]), .Ci(1'b0) );
endmodule


module ADDER_P4_N_BIT64_2 ( A, B, add_sub, Cout, SUM );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input add_sub;
  output Cout;

  wire   [63:0] B_xor;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31;
  assign B_xor[31] = B[31];
  assign B_xor[30] = B[30];
  assign B_xor[29] = B[29];
  assign B_xor[28] = B[28];
  assign B_xor[27] = B[27];
  assign B_xor[26] = B[26];
  assign B_xor[25] = B[25];
  assign B_xor[24] = B[24];
  assign B_xor[23] = B[23];
  assign B_xor[22] = B[22];
  assign B_xor[21] = B[21];
  assign B_xor[20] = B[20];
  assign B_xor[19] = B[19];
  assign B_xor[18] = B[18];
  assign B_xor[17] = B[17];
  assign B_xor[16] = B[16];
  assign B_xor[15] = B[15];
  assign B_xor[14] = B[14];
  assign B_xor[13] = B[13];
  assign B_xor[12] = B[12];
  assign B_xor[11] = B[11];
  assign B_xor[10] = B[10];
  assign B_xor[9] = B[9];
  assign B_xor[8] = B[8];
  assign B_xor[7] = B[7];
  assign B_xor[6] = B[6];
  assign B_xor[5] = B[5];
  assign B_xor[4] = B[4];
  assign B_xor[3] = B[3];
  assign B_xor[2] = B[2];
  assign B_xor[1] = B[1];
  assign B_xor[0] = B[0];

  SUMGENERATOR_Nblocks16_bits_per_block4_2 CSA ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, A[31:28], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B_xor[31:0]}), 
        .CARRY_SELECT({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .SUM({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, SUM[31:0]}) );
endmodule


module FA_128 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_127 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_126 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_125 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_32 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_128 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_127 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_126 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_125 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_16 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_16 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_32 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0) );
  MUX_2to1_N4_16 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_120 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_119 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_118 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_117 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_30 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_120 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_119 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_118 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_117 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_15 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_15 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_30 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0) );
  MUX_2to1_N4_15 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_112 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_111 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_110 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_109 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_28 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_112 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_111 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_110 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_109 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_14 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_14 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_28 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0) );
  MUX_2to1_N4_14 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_104 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_103 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_102 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_101 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_26 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_104 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_103 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_102 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_101 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_13 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_13 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_26 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0) );
  MUX_2to1_N4_13 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_96 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_95 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_94 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_93 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_24 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_96 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_95 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_94 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_93 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_12 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_12 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_24 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0) );
  MUX_2to1_N4_12 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_88 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_87 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_86 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_85 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_22 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_88 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_87 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_86 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_85 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_11 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_11 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_22 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0) );
  MUX_2to1_N4_11 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_80 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_79 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_78 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_77 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module RCA_N4_20 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;


  FA_80 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_79 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_78 FULLADDER_3 ( .A(1'b0), .B(B[2]), .Ci(1'b0), .S(S[2]) );
  FA_77 FULLADDER_4 ( .A(1'b0), .B(B[3]), .Ci(1'b0), .S(S[3]) );
endmodule


module MUX_2to1_N4_10 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_10 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_20 RCA_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0) );
  MUX_2to1_N4_10 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module FA_72 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_71 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   B;
  assign S = B;

endmodule


module FA_70 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(S) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(Co) );
endmodule


module FA_69 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n1;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n1) );
  XNOR2_X1 U2 ( .A(n1), .B(Ci), .ZN(S) );
endmodule


module RCA_N4_18 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;
  wire   \CTMP[3] ;

  FA_72 FULLADDER_1 ( .A(1'b0), .B(B[0]), .Ci(1'b0), .S(S[0]) );
  FA_71 FULLADDER_2 ( .A(1'b0), .B(B[1]), .Ci(1'b0), .S(S[1]) );
  FA_70 FULLADDER_3 ( .A(A[2]), .B(B[2]), .Ci(1'b0), .S(S[2]), .Co(\CTMP[3] )
         );
  FA_69 FULLADDER_4 ( .A(A[3]), .B(B[3]), .Ci(\CTMP[3] ), .S(S[3]) );
endmodule


module MUX_2to1_N4_9 ( IN0, IN1, SEL, Y );
  input [3:0] IN0;
  input [3:0] IN1;
  output [3:0] Y;
  input SEL;

  assign Y[3] = IN0[3];
  assign Y[2] = IN0[2];
  assign Y[1] = IN0[1];
  assign Y[0] = IN0[0];

endmodule


module carry_select_block_N4_9 ( A, B, S, Ci );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S_0;

  RCA_N4_18 RCA_0 ( .A({A[3:2], 1'b0, 1'b0}), .B(B), .Ci(1'b0), .S(S_0) );
  MUX_2to1_N4_9 SUM_SELECT_MUX ( .IN0(S_0), .IN1({1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(1'b0), .Y(S) );
endmodule


module SUMGENERATOR_Nblocks16_bits_per_block4_1 ( A, B, CARRY_SELECT, SUM );
  input [63:0] A;
  input [63:0] B;
  input [15:0] CARRY_SELECT;
  output [63:0] SUM;


  carry_select_block_N4_16 block_n_1 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B[3:0]), .S(SUM[3:0]), .Ci(1'b0) );
  carry_select_block_N4_15 block_n_2 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(B[7:4]), .S(SUM[7:4]), .Ci(1'b0) );
  carry_select_block_N4_14 block_n_3 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(
        B[11:8]), .S(SUM[11:8]), .Ci(1'b0) );
  carry_select_block_N4_13 block_n_4 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(
        B[15:12]), .S(SUM[15:12]), .Ci(1'b0) );
  carry_select_block_N4_12 block_n_5 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(
        B[19:16]), .S(SUM[19:16]), .Ci(1'b0) );
  carry_select_block_N4_11 block_n_6 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(
        B[23:20]), .S(SUM[23:20]), .Ci(1'b0) );
  carry_select_block_N4_10 block_n_7 ( .A({1'b0, 1'b0, 1'b0, 1'b0}), .B(
        B[27:24]), .S(SUM[27:24]), .Ci(1'b0) );
  carry_select_block_N4_9 block_n_8 ( .A({A[31:30], 1'b0, 1'b0}), .B(B[31:28]), 
        .S(SUM[31:28]), .Ci(1'b0) );
endmodule


module ADDER_P4_N_BIT64_1 ( A, B, add_sub, Cout, SUM );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input add_sub;
  output Cout;

  wire   [63:0] B_xor;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31;
  assign B_xor[31] = B[31];
  assign B_xor[30] = B[30];
  assign B_xor[29] = B[29];
  assign B_xor[28] = B[28];
  assign B_xor[27] = B[27];
  assign B_xor[26] = B[26];
  assign B_xor[25] = B[25];
  assign B_xor[24] = B[24];
  assign B_xor[23] = B[23];
  assign B_xor[22] = B[22];
  assign B_xor[21] = B[21];
  assign B_xor[20] = B[20];
  assign B_xor[19] = B[19];
  assign B_xor[18] = B[18];
  assign B_xor[17] = B[17];
  assign B_xor[16] = B[16];
  assign B_xor[15] = B[15];
  assign B_xor[14] = B[14];
  assign B_xor[13] = B[13];
  assign B_xor[12] = B[12];
  assign B_xor[11] = B[11];
  assign B_xor[10] = B[10];
  assign B_xor[9] = B[9];
  assign B_xor[8] = B[8];
  assign B_xor[7] = B[7];
  assign B_xor[6] = B[6];
  assign B_xor[5] = B[5];
  assign B_xor[4] = B[4];
  assign B_xor[3] = B[3];
  assign B_xor[2] = B[2];
  assign B_xor[1] = B[1];
  assign B_xor[0] = B[0];

  SUMGENERATOR_Nblocks16_bits_per_block4_1 CSA ( .A({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, A[31:30], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, B_xor[31:0]}), 
        .CARRY_SELECT({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .SUM({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, SUM[31:0]}) );
endmodule


module MUX_8to1_N64_0 ( IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, SEL, Y );
  input [63:0] IN0;
  input [63:0] IN1;
  input [63:0] IN2;
  input [63:0] IN3;
  input [63:0] IN4;
  input [63:0] IN5;
  input [63:0] IN6;
  input [63:0] IN7;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107;

  BUF_X2 U1 ( .A(n105), .Z(n50) );
  NAND2_X1 U2 ( .A1(n54), .A2(n53), .ZN(Y[10]) );
  BUF_X1 U3 ( .A(n103), .Z(n14) );
  INV_X1 U4 ( .A(n12), .ZN(n13) );
  AOI22_X1 U5 ( .A1(n49), .A2(IN1[17]), .B1(IN4[18]), .B2(n50), .ZN(n1) );
  AOI22_X1 U6 ( .A1(IN4[19]), .A2(n47), .B1(n46), .B2(IN1[18]), .ZN(n2) );
  NAND2_X1 U7 ( .A1(n1), .A2(n2), .ZN(Y[18]) );
  AOI22_X1 U8 ( .A1(n49), .A2(IN1[18]), .B1(n50), .B2(IN4[19]), .ZN(n3) );
  AOI22_X1 U9 ( .A1(IN4[20]), .A2(n47), .B1(n46), .B2(IN1[19]), .ZN(n4) );
  NAND2_X1 U10 ( .A1(n3), .A2(n4), .ZN(Y[19]) );
  AOI22_X1 U11 ( .A1(n49), .A2(IN1[22]), .B1(IN4[23]), .B2(n50), .ZN(n5) );
  AOI22_X1 U12 ( .A1(IN4[24]), .A2(n47), .B1(n46), .B2(IN1[23]), .ZN(n6) );
  NAND2_X1 U13 ( .A1(n5), .A2(n6), .ZN(Y[23]) );
  AOI22_X1 U14 ( .A1(n49), .A2(IN1[12]), .B1(n50), .B2(IN4[13]), .ZN(n7) );
  AOI22_X1 U15 ( .A1(IN4[14]), .A2(n47), .B1(n46), .B2(IN1[13]), .ZN(n8) );
  NAND2_X1 U16 ( .A1(n7), .A2(n8), .ZN(Y[13]) );
  NAND2_X1 U17 ( .A1(IN4[6]), .A2(n103), .ZN(n9) );
  NAND2_X1 U18 ( .A1(IN1[5]), .A2(n45), .ZN(n10) );
  NAND3_X1 U19 ( .A1(n10), .A2(n96), .A3(n9), .ZN(Y[5]) );
  BUF_X1 U20 ( .A(n48), .Z(n11) );
  CLKBUF_X1 U21 ( .A(n48), .Z(n32) );
  AND3_X1 U22 ( .A1(SEL[2]), .A2(n36), .A3(n52), .ZN(n105) );
  INV_X1 U23 ( .A(n50), .ZN(n12) );
  BUF_X2 U24 ( .A(n102), .Z(n45) );
  CLKBUF_X3 U25 ( .A(n102), .Z(n46) );
  NAND2_X1 U26 ( .A1(n63), .A2(n62), .ZN(Y[16]) );
  AND2_X1 U27 ( .A1(n46), .A2(IN1[25]), .ZN(n37) );
  INV_X1 U28 ( .A(SEL[0]), .ZN(n52) );
  NAND2_X1 U29 ( .A1(n101), .A2(n30), .ZN(Y[8]) );
  AOI22_X1 U30 ( .A1(n47), .A2(IN4[9]), .B1(n46), .B2(IN1[8]), .ZN(n30) );
  BUF_X1 U31 ( .A(n49), .Z(n31) );
  AND2_X1 U32 ( .A1(SEL[1]), .A2(n33), .ZN(n103) );
  INV_X1 U33 ( .A(SEL[1]), .ZN(n36) );
  NOR2_X1 U34 ( .A1(SEL[0]), .A2(SEL[2]), .ZN(n33) );
  NOR2_X1 U35 ( .A1(n34), .A2(n52), .ZN(n104) );
  NAND2_X1 U36 ( .A1(n35), .A2(SEL[1]), .ZN(n34) );
  INV_X1 U37 ( .A(SEL[2]), .ZN(n35) );
  AOI21_X1 U38 ( .B1(IN4[26]), .B2(n47), .A(n37), .ZN(n77) );
  BUF_X4 U39 ( .A(n103), .Z(n47) );
  BUF_X2 U40 ( .A(n104), .Z(n48) );
  BUF_X2 U41 ( .A(n104), .Z(n49) );
  AND2_X1 U42 ( .A1(n46), .A2(IN1[10]), .ZN(n38) );
  AOI21_X1 U43 ( .B1(IN4[11]), .B2(n47), .A(n38), .ZN(n54) );
  NAND2_X1 U44 ( .A1(n55), .A2(n39), .ZN(Y[11]) );
  AOI21_X1 U45 ( .B1(IN4[12]), .B2(n47), .A(n40), .ZN(n39) );
  AND2_X1 U46 ( .A1(n46), .A2(IN1[11]), .ZN(n40) );
  AOI21_X1 U47 ( .B1(IN4[21]), .B2(n47), .A(n41), .ZN(n69) );
  AND2_X1 U48 ( .A1(n46), .A2(IN1[20]), .ZN(n41) );
  AOI21_X1 U49 ( .B1(IN4[23]), .B2(n47), .A(n42), .ZN(n73) );
  AND2_X1 U50 ( .A1(n46), .A2(IN1[22]), .ZN(n42) );
  AOI21_X1 U51 ( .B1(IN4[22]), .B2(n47), .A(n43), .ZN(n71) );
  AND2_X1 U52 ( .A1(n46), .A2(IN1[21]), .ZN(n43) );
  AOI21_X1 U53 ( .B1(IN4[16]), .B2(n47), .A(n44), .ZN(n61) );
  AND2_X1 U54 ( .A1(n46), .A2(IN1[15]), .ZN(n44) );
  NOR3_X1 U55 ( .A1(n52), .A2(SEL[2]), .A3(SEL[1]), .ZN(n102) );
  OAI21_X1 U56 ( .B1(n46), .B2(n47), .A(IN1[0]), .ZN(n51) );
  INV_X1 U57 ( .A(n51), .ZN(Y[0]) );
  AOI22_X1 U58 ( .A1(n50), .A2(IN4[10]), .B1(n32), .B2(IN1[9]), .ZN(n53) );
  AOI22_X1 U59 ( .A1(n50), .A2(IN4[11]), .B1(n49), .B2(IN1[10]), .ZN(n55) );
  AOI22_X1 U60 ( .A1(n46), .A2(IN1[12]), .B1(IN4[13]), .B2(n47), .ZN(n57) );
  AOI22_X1 U61 ( .A1(IN4[12]), .A2(n50), .B1(n49), .B2(IN1[11]), .ZN(n56) );
  NAND2_X1 U62 ( .A1(n56), .A2(n57), .ZN(Y[12]) );
  AOI22_X1 U63 ( .A1(n46), .A2(IN1[14]), .B1(n47), .B2(IN4[15]), .ZN(n59) );
  AOI22_X1 U64 ( .A1(n50), .A2(IN4[14]), .B1(n49), .B2(IN1[13]), .ZN(n58) );
  NAND2_X1 U65 ( .A1(n59), .A2(n58), .ZN(Y[14]) );
  AOI22_X1 U66 ( .A1(n50), .A2(IN4[15]), .B1(n49), .B2(IN1[14]), .ZN(n60) );
  NAND2_X1 U67 ( .A1(n61), .A2(n60), .ZN(Y[15]) );
  AOI22_X1 U68 ( .A1(n46), .A2(IN1[16]), .B1(n47), .B2(IN4[17]), .ZN(n63) );
  AOI22_X1 U69 ( .A1(IN4[16]), .A2(n50), .B1(n49), .B2(IN1[15]), .ZN(n62) );
  AOI22_X1 U70 ( .A1(n46), .A2(IN1[17]), .B1(n47), .B2(IN4[18]), .ZN(n65) );
  AOI22_X1 U71 ( .A1(n50), .A2(IN4[17]), .B1(n49), .B2(IN1[16]), .ZN(n64) );
  NAND2_X1 U72 ( .A1(n65), .A2(n64), .ZN(Y[17]) );
  OAI21_X1 U73 ( .B1(n13), .B2(n31), .A(IN1[0]), .ZN(n67) );
  AOI22_X1 U74 ( .A1(n46), .A2(IN1[1]), .B1(n47), .B2(IN4[2]), .ZN(n66) );
  NAND2_X1 U75 ( .A1(n67), .A2(n66), .ZN(Y[1]) );
  AOI22_X1 U76 ( .A1(IN4[20]), .A2(n50), .B1(n49), .B2(IN1[19]), .ZN(n68) );
  NAND2_X1 U77 ( .A1(n69), .A2(n68), .ZN(Y[20]) );
  AOI22_X1 U78 ( .A1(IN4[21]), .A2(n50), .B1(n49), .B2(IN1[20]), .ZN(n70) );
  NAND2_X1 U79 ( .A1(n71), .A2(n70), .ZN(Y[21]) );
  AOI22_X1 U80 ( .A1(n50), .A2(IN4[22]), .B1(n49), .B2(IN1[21]), .ZN(n72) );
  NAND2_X1 U81 ( .A1(n73), .A2(n72), .ZN(Y[22]) );
  AOI22_X1 U82 ( .A1(n46), .A2(IN1[24]), .B1(n47), .B2(IN4[25]), .ZN(n75) );
  AOI22_X1 U83 ( .A1(n13), .A2(IN4[24]), .B1(n49), .B2(IN1[23]), .ZN(n74) );
  NAND2_X1 U84 ( .A1(n75), .A2(n74), .ZN(Y[24]) );
  AOI22_X1 U85 ( .A1(IN4[25]), .A2(n13), .B1(n49), .B2(IN1[24]), .ZN(n76) );
  NAND2_X1 U86 ( .A1(n77), .A2(n76), .ZN(Y[25]) );
  AOI22_X1 U87 ( .A1(n46), .A2(IN1[26]), .B1(n47), .B2(IN4[27]), .ZN(n79) );
  AOI22_X1 U88 ( .A1(IN4[26]), .A2(n13), .B1(n31), .B2(IN1[25]), .ZN(n78) );
  NAND2_X1 U89 ( .A1(n79), .A2(n78), .ZN(Y[26]) );
  AOI22_X1 U90 ( .A1(n46), .A2(IN1[27]), .B1(IN4[28]), .B2(n47), .ZN(n81) );
  AOI22_X1 U91 ( .A1(n13), .A2(IN4[27]), .B1(n31), .B2(IN1[26]), .ZN(n80) );
  NAND2_X1 U92 ( .A1(n81), .A2(n80), .ZN(Y[27]) );
  AOI22_X1 U93 ( .A1(n46), .A2(IN1[28]), .B1(n47), .B2(IN4[29]), .ZN(n83) );
  AOI22_X1 U94 ( .A1(IN4[28]), .A2(n13), .B1(n31), .B2(IN1[27]), .ZN(n82) );
  NAND2_X1 U95 ( .A1(n83), .A2(n82), .ZN(Y[28]) );
  AOI22_X1 U96 ( .A1(n45), .A2(IN1[29]), .B1(n47), .B2(IN4[30]), .ZN(n85) );
  AOI22_X1 U97 ( .A1(n13), .A2(IN4[29]), .B1(n32), .B2(IN1[28]), .ZN(n84) );
  NAND2_X1 U98 ( .A1(n85), .A2(n84), .ZN(Y[29]) );
  AOI22_X1 U99 ( .A1(n46), .A2(IN1[2]), .B1(n47), .B2(IN4[3]), .ZN(n87) );
  AOI22_X1 U100 ( .A1(n50), .A2(IN4[2]), .B1(n32), .B2(IN1[1]), .ZN(n86) );
  NAND2_X1 U101 ( .A1(n87), .A2(n86), .ZN(Y[2]) );
  AOI22_X1 U102 ( .A1(n46), .A2(IN1[30]), .B1(n47), .B2(IN4[31]), .ZN(n89) );
  AOI22_X1 U103 ( .A1(n13), .A2(IN4[30]), .B1(n32), .B2(IN1[29]), .ZN(n88) );
  NAND2_X1 U104 ( .A1(n89), .A2(n88), .ZN(Y[30]) );
  AOI22_X1 U105 ( .A1(n46), .A2(IN1[31]), .B1(n47), .B2(IN2[31]), .ZN(n91) );
  AOI22_X1 U106 ( .A1(n13), .A2(IN4[31]), .B1(n32), .B2(IN1[30]), .ZN(n90) );
  NAND2_X1 U107 ( .A1(n91), .A2(n90), .ZN(Y[31]) );
  AOI22_X1 U108 ( .A1(n45), .A2(IN1[3]), .B1(n14), .B2(IN4[4]), .ZN(n93) );
  AOI22_X1 U109 ( .A1(n105), .A2(IN4[3]), .B1(n11), .B2(IN1[2]), .ZN(n92) );
  NAND2_X1 U110 ( .A1(n93), .A2(n92), .ZN(Y[3]) );
  AOI22_X1 U111 ( .A1(n45), .A2(IN1[4]), .B1(n14), .B2(IN4[5]), .ZN(n95) );
  AOI22_X1 U112 ( .A1(n105), .A2(IN4[4]), .B1(n48), .B2(IN1[3]), .ZN(n94) );
  NAND2_X1 U113 ( .A1(n95), .A2(n94), .ZN(Y[4]) );
  AOI22_X1 U114 ( .A1(n105), .A2(IN4[5]), .B1(n104), .B2(IN1[4]), .ZN(n96) );
  AOI22_X1 U115 ( .A1(n45), .A2(IN1[6]), .B1(n14), .B2(IN4[7]), .ZN(n98) );
  AOI22_X1 U116 ( .A1(n105), .A2(IN4[6]), .B1(n48), .B2(IN1[5]), .ZN(n97) );
  NAND2_X1 U117 ( .A1(n98), .A2(n97), .ZN(Y[6]) );
  AOI22_X1 U118 ( .A1(n45), .A2(IN1[7]), .B1(n14), .B2(IN4[8]), .ZN(n100) );
  AOI22_X1 U119 ( .A1(n105), .A2(IN4[7]), .B1(n48), .B2(IN1[6]), .ZN(n99) );
  NAND2_X1 U120 ( .A1(n99), .A2(n100), .ZN(Y[7]) );
  AOI22_X1 U121 ( .A1(n105), .A2(IN4[8]), .B1(n49), .B2(IN1[7]), .ZN(n101) );
  AOI22_X1 U122 ( .A1(n47), .A2(IN4[10]), .B1(IN1[9]), .B2(n46), .ZN(n107) );
  AOI22_X1 U123 ( .A1(n50), .A2(IN4[9]), .B1(n49), .B2(IN1[8]), .ZN(n106) );
  NAND2_X1 U124 ( .A1(n107), .A2(n106), .ZN(Y[9]) );
endmodule


module MUX_8to1_N64_15 ( IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, SEL, Y );
  input [63:0] IN0;
  input [63:0] IN1;
  input [63:0] IN2;
  input [63:0] IN3;
  input [63:0] IN4;
  input [63:0] IN5;
  input [63:0] IN6;
  input [63:0] IN7;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n1, n2, n3, n4, n5, n6, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97;

  BUF_X1 U1 ( .A(n92), .Z(n1) );
  BUF_X1 U2 ( .A(n92), .Z(n2) );
  AND3_X2 U3 ( .A1(n23), .A2(n24), .A3(SEL[0]), .ZN(n92) );
  BUF_X1 U4 ( .A(n92), .Z(n29) );
  BUF_X4 U5 ( .A(n28), .Z(n27) );
  BUF_X1 U6 ( .A(n95), .Z(n35) );
  BUF_X2 U7 ( .A(n93), .Z(n32) );
  AOI22_X1 U8 ( .A1(n34), .A2(IN1[14]), .B1(IN4[15]), .B2(n36), .ZN(n3) );
  AOI22_X1 U9 ( .A1(IN4[16]), .A2(n31), .B1(n29), .B2(IN1[15]), .ZN(n4) );
  NAND2_X1 U10 ( .A1(n3), .A2(n4), .ZN(Y[15]) );
  AOI22_X1 U11 ( .A1(n92), .A2(IN1[3]), .B1(n32), .B2(IN4[4]), .ZN(n5) );
  OAI21_X1 U12 ( .B1(n37), .B2(n33), .A(IN1[2]), .ZN(n6) );
  NAND2_X1 U13 ( .A1(n6), .A2(n5), .ZN(Y[3]) );
  BUF_X4 U14 ( .A(n94), .Z(n34) );
  CLKBUF_X3 U15 ( .A(n95), .Z(n36) );
  NAND2_X1 U16 ( .A1(n40), .A2(n41), .ZN(Y[4]) );
  BUF_X1 U17 ( .A(n35), .Z(n22) );
  NAND2_X1 U18 ( .A1(n42), .A2(n43), .ZN(Y[5]) );
  NAND2_X1 U19 ( .A1(n46), .A2(n47), .ZN(Y[7]) );
  OR2_X1 U20 ( .A1(SEL[0]), .A2(SEL[2]), .ZN(n25) );
  INV_X1 U21 ( .A(SEL[1]), .ZN(n23) );
  INV_X1 U22 ( .A(SEL[2]), .ZN(n24) );
  BUF_X2 U23 ( .A(n94), .Z(n33) );
  AND3_X1 U24 ( .A1(n24), .A2(SEL[1]), .A3(SEL[0]), .ZN(n94) );
  NOR2_X1 U25 ( .A1(n25), .A2(n23), .ZN(n93) );
  CLKBUF_X3 U26 ( .A(n93), .Z(n31) );
  BUF_X2 U27 ( .A(n92), .Z(n28) );
  BUF_X2 U28 ( .A(n95), .Z(n37) );
  BUF_X1 U29 ( .A(n31), .Z(n30) );
  AOI21_X1 U30 ( .B1(IN4[13]), .B2(n31), .A(n26), .ZN(n57) );
  AND2_X1 U31 ( .A1(n92), .A2(IN1[12]), .ZN(n26) );
  INV_X1 U32 ( .A(SEL[0]), .ZN(n39) );
  OAI21_X1 U33 ( .B1(n28), .B2(n31), .A(IN1[2]), .ZN(n38) );
  INV_X1 U34 ( .A(n38), .ZN(Y[2]) );
  AND3_X1 U35 ( .A1(n23), .A2(SEL[2]), .A3(n39), .ZN(n95) );
  AOI22_X1 U36 ( .A1(n32), .A2(IN4[5]), .B1(n92), .B2(IN1[4]), .ZN(n41) );
  AOI22_X1 U37 ( .A1(IN4[4]), .A2(n37), .B1(n33), .B2(IN1[3]), .ZN(n40) );
  AOI22_X1 U38 ( .A1(n32), .A2(IN4[6]), .B1(n92), .B2(IN1[5]), .ZN(n43) );
  AOI22_X1 U39 ( .A1(n95), .A2(IN4[5]), .B1(n33), .B2(IN1[4]), .ZN(n42) );
  AOI22_X1 U40 ( .A1(n32), .A2(IN4[7]), .B1(n92), .B2(IN1[6]), .ZN(n45) );
  AOI22_X1 U41 ( .A1(n37), .A2(IN4[6]), .B1(n33), .B2(IN1[5]), .ZN(n44) );
  NAND2_X1 U42 ( .A1(n45), .A2(n44), .ZN(Y[6]) );
  AOI22_X1 U43 ( .A1(n32), .A2(IN4[8]), .B1(n92), .B2(IN1[7]), .ZN(n47) );
  AOI22_X1 U44 ( .A1(n37), .A2(IN4[7]), .B1(n33), .B2(IN1[6]), .ZN(n46) );
  AOI22_X1 U45 ( .A1(n31), .A2(IN4[9]), .B1(n92), .B2(IN1[8]), .ZN(n49) );
  AOI22_X1 U46 ( .A1(n35), .A2(IN4[8]), .B1(n33), .B2(IN1[7]), .ZN(n48) );
  NAND2_X1 U47 ( .A1(n49), .A2(n48), .ZN(Y[8]) );
  AOI22_X1 U48 ( .A1(n32), .A2(IN4[10]), .B1(n92), .B2(IN1[9]), .ZN(n51) );
  AOI22_X1 U49 ( .A1(n37), .A2(IN4[9]), .B1(n33), .B2(IN1[8]), .ZN(n50) );
  NAND2_X1 U50 ( .A1(n51), .A2(n50), .ZN(Y[9]) );
  AOI22_X1 U51 ( .A1(n31), .A2(IN4[11]), .B1(n92), .B2(IN1[10]), .ZN(n53) );
  AOI22_X1 U52 ( .A1(n35), .A2(IN4[10]), .B1(n34), .B2(IN1[9]), .ZN(n52) );
  NAND2_X1 U53 ( .A1(n53), .A2(n52), .ZN(Y[10]) );
  AOI22_X1 U54 ( .A1(n31), .A2(IN4[12]), .B1(n92), .B2(IN1[11]), .ZN(n55) );
  AOI22_X1 U55 ( .A1(n36), .A2(IN4[11]), .B1(n34), .B2(IN1[10]), .ZN(n54) );
  NAND2_X1 U56 ( .A1(n55), .A2(n54), .ZN(Y[11]) );
  AOI22_X1 U57 ( .A1(IN4[12]), .A2(n36), .B1(n34), .B2(IN1[11]), .ZN(n56) );
  NAND2_X1 U58 ( .A1(n57), .A2(n56), .ZN(Y[12]) );
  AOI22_X1 U59 ( .A1(IN4[14]), .A2(n31), .B1(n1), .B2(IN1[13]), .ZN(n59) );
  AOI22_X1 U60 ( .A1(n36), .A2(IN4[13]), .B1(n34), .B2(IN1[12]), .ZN(n58) );
  NAND2_X1 U61 ( .A1(n59), .A2(n58), .ZN(Y[13]) );
  AOI22_X1 U62 ( .A1(n31), .A2(IN4[15]), .B1(n2), .B2(IN1[14]), .ZN(n61) );
  AOI22_X1 U63 ( .A1(n36), .A2(IN4[14]), .B1(n34), .B2(IN1[13]), .ZN(n60) );
  NAND2_X1 U64 ( .A1(n61), .A2(n60), .ZN(Y[14]) );
  AOI22_X1 U65 ( .A1(n31), .A2(IN4[17]), .B1(n28), .B2(IN1[16]), .ZN(n63) );
  AOI22_X1 U66 ( .A1(n36), .A2(IN4[16]), .B1(n34), .B2(IN1[15]), .ZN(n62) );
  NAND2_X1 U67 ( .A1(n63), .A2(n62), .ZN(Y[16]) );
  AOI22_X1 U68 ( .A1(n31), .A2(IN4[18]), .B1(n28), .B2(IN1[17]), .ZN(n65) );
  AOI22_X1 U69 ( .A1(n35), .A2(IN4[17]), .B1(n34), .B2(IN1[16]), .ZN(n64) );
  NAND2_X1 U70 ( .A1(n65), .A2(n64), .ZN(Y[17]) );
  AOI22_X1 U71 ( .A1(n31), .A2(IN4[19]), .B1(n28), .B2(IN1[18]), .ZN(n67) );
  AOI22_X1 U72 ( .A1(n36), .A2(IN4[18]), .B1(n34), .B2(IN1[17]), .ZN(n66) );
  NAND2_X1 U73 ( .A1(n67), .A2(n66), .ZN(Y[18]) );
  AOI22_X1 U74 ( .A1(n31), .A2(IN4[20]), .B1(n28), .B2(IN1[19]), .ZN(n69) );
  AOI22_X1 U75 ( .A1(n36), .A2(IN4[19]), .B1(n34), .B2(IN1[18]), .ZN(n68) );
  NAND2_X1 U76 ( .A1(n69), .A2(n68), .ZN(Y[19]) );
  AOI22_X1 U77 ( .A1(n31), .A2(IN4[21]), .B1(n28), .B2(IN1[20]), .ZN(n71) );
  AOI22_X1 U78 ( .A1(n36), .A2(IN4[20]), .B1(n34), .B2(IN1[19]), .ZN(n70) );
  NAND2_X1 U79 ( .A1(n71), .A2(n70), .ZN(Y[20]) );
  AOI22_X1 U80 ( .A1(n30), .A2(IN4[22]), .B1(n1), .B2(IN1[21]), .ZN(n73) );
  AOI22_X1 U81 ( .A1(n35), .A2(IN4[21]), .B1(n34), .B2(IN1[20]), .ZN(n72) );
  NAND2_X1 U82 ( .A1(n73), .A2(n72), .ZN(Y[21]) );
  AOI22_X1 U83 ( .A1(n30), .A2(IN4[23]), .B1(n27), .B2(IN1[22]), .ZN(n75) );
  AOI22_X1 U84 ( .A1(n35), .A2(IN4[22]), .B1(n34), .B2(IN1[21]), .ZN(n74) );
  NAND2_X1 U85 ( .A1(n75), .A2(n74), .ZN(Y[22]) );
  AOI22_X1 U86 ( .A1(n30), .A2(IN4[24]), .B1(n27), .B2(IN1[23]), .ZN(n77) );
  AOI22_X1 U87 ( .A1(n35), .A2(IN4[23]), .B1(n34), .B2(IN1[22]), .ZN(n76) );
  NAND2_X1 U88 ( .A1(n77), .A2(n76), .ZN(Y[23]) );
  AOI22_X1 U89 ( .A1(n30), .A2(IN4[25]), .B1(n27), .B2(IN1[24]), .ZN(n79) );
  AOI22_X1 U90 ( .A1(IN4[24]), .A2(n22), .B1(n34), .B2(IN1[23]), .ZN(n78) );
  NAND2_X1 U91 ( .A1(n79), .A2(n78), .ZN(Y[24]) );
  AOI22_X1 U92 ( .A1(n30), .A2(IN4[26]), .B1(n27), .B2(IN1[25]), .ZN(n81) );
  AOI22_X1 U93 ( .A1(n22), .A2(IN4[25]), .B1(n34), .B2(IN1[24]), .ZN(n80) );
  NAND2_X1 U94 ( .A1(n81), .A2(n80), .ZN(Y[25]) );
  AOI22_X1 U95 ( .A1(n30), .A2(IN4[27]), .B1(n27), .B2(IN1[26]), .ZN(n83) );
  AOI22_X1 U96 ( .A1(n22), .A2(IN4[26]), .B1(n34), .B2(IN1[25]), .ZN(n82) );
  NAND2_X1 U97 ( .A1(n83), .A2(n82), .ZN(Y[26]) );
  AOI22_X1 U98 ( .A1(n30), .A2(IN4[28]), .B1(n27), .B2(IN1[27]), .ZN(n85) );
  AOI22_X1 U99 ( .A1(n22), .A2(IN4[27]), .B1(n34), .B2(IN1[26]), .ZN(n84) );
  NAND2_X1 U100 ( .A1(n85), .A2(n84), .ZN(Y[27]) );
  AOI22_X1 U101 ( .A1(n30), .A2(IN4[29]), .B1(n27), .B2(IN1[28]), .ZN(n87) );
  AOI22_X1 U102 ( .A1(n22), .A2(IN4[28]), .B1(n34), .B2(IN1[27]), .ZN(n86) );
  NAND2_X1 U103 ( .A1(n87), .A2(n86), .ZN(Y[28]) );
  AOI22_X1 U104 ( .A1(n30), .A2(IN4[30]), .B1(n27), .B2(IN1[29]), .ZN(n89) );
  AOI22_X1 U105 ( .A1(n22), .A2(IN4[29]), .B1(n34), .B2(IN1[28]), .ZN(n88) );
  NAND2_X1 U106 ( .A1(n89), .A2(n88), .ZN(Y[29]) );
  AOI22_X1 U107 ( .A1(n30), .A2(IN4[31]), .B1(n27), .B2(IN1[30]), .ZN(n91) );
  AOI22_X1 U108 ( .A1(n22), .A2(IN4[30]), .B1(n34), .B2(IN1[29]), .ZN(n90) );
  NAND2_X1 U109 ( .A1(n91), .A2(n90), .ZN(Y[30]) );
  AOI22_X1 U110 ( .A1(n30), .A2(IN2[31]), .B1(n27), .B2(IN1[31]), .ZN(n97) );
  AOI22_X1 U111 ( .A1(n36), .A2(IN4[31]), .B1(n34), .B2(IN1[30]), .ZN(n96) );
  NAND2_X1 U112 ( .A1(n97), .A2(n96), .ZN(Y[31]) );
endmodule


module MUX_8to1_N64_14 ( IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, SEL, Y );
  input [63:0] IN0;
  input [63:0] IN1;
  input [63:0] IN2;
  input [63:0] IN3;
  input [63:0] IN4;
  input [63:0] IN5;
  input [63:0] IN6;
  input [63:0] IN7;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n12, n14, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82;

  NAND2_X1 U1 ( .A1(n68), .A2(n67), .ZN(Y[26]) );
  BUF_X2 U2 ( .A(n79), .Z(n12) );
  BUF_X2 U3 ( .A(n78), .Z(n14) );
  AND3_X2 U4 ( .A1(n24), .A2(n23), .A3(SEL[2]), .ZN(n80) );
  BUF_X1 U5 ( .A(n77), .Z(n21) );
  NOR3_X1 U6 ( .A1(SEL[2]), .A2(SEL[1]), .A3(n23), .ZN(n77) );
  INV_X1 U7 ( .A(SEL[1]), .ZN(n24) );
  NOR3_X1 U8 ( .A1(SEL[2]), .A2(SEL[0]), .A3(n24), .ZN(n78) );
  INV_X1 U9 ( .A(SEL[0]), .ZN(n23) );
  OAI21_X1 U10 ( .B1(n14), .B2(n77), .A(IN1[4]), .ZN(n22) );
  INV_X1 U11 ( .A(n22), .ZN(Y[4]) );
  NOR3_X1 U12 ( .A1(SEL[2]), .A2(n24), .A3(n23), .ZN(n79) );
  OAI21_X1 U13 ( .B1(n80), .B2(n12), .A(IN1[4]), .ZN(n26) );
  AOI22_X1 U14 ( .A1(n14), .A2(IN4[6]), .B1(n21), .B2(IN1[5]), .ZN(n25) );
  NAND2_X1 U15 ( .A1(n26), .A2(n25), .ZN(Y[5]) );
  AOI22_X1 U16 ( .A1(n14), .A2(IN4[7]), .B1(n77), .B2(IN1[6]), .ZN(n28) );
  AOI22_X1 U17 ( .A1(IN4[6]), .A2(n80), .B1(n12), .B2(IN1[5]), .ZN(n27) );
  NAND2_X1 U18 ( .A1(n28), .A2(n27), .ZN(Y[6]) );
  AOI22_X1 U19 ( .A1(n14), .A2(IN4[8]), .B1(n77), .B2(IN1[7]), .ZN(n30) );
  AOI22_X1 U20 ( .A1(n80), .A2(IN4[7]), .B1(n12), .B2(IN1[6]), .ZN(n29) );
  NAND2_X1 U21 ( .A1(n30), .A2(n29), .ZN(Y[7]) );
  AOI22_X1 U22 ( .A1(n14), .A2(IN4[9]), .B1(n77), .B2(IN1[8]), .ZN(n32) );
  AOI22_X1 U23 ( .A1(n80), .A2(IN4[8]), .B1(n12), .B2(IN1[7]), .ZN(n31) );
  NAND2_X1 U24 ( .A1(n32), .A2(n31), .ZN(Y[8]) );
  AOI22_X1 U25 ( .A1(n14), .A2(IN4[10]), .B1(n21), .B2(IN1[9]), .ZN(n34) );
  AOI22_X1 U26 ( .A1(n80), .A2(IN4[9]), .B1(n12), .B2(IN1[8]), .ZN(n33) );
  NAND2_X1 U27 ( .A1(n34), .A2(n33), .ZN(Y[9]) );
  AOI22_X1 U28 ( .A1(n14), .A2(IN4[11]), .B1(n21), .B2(IN1[10]), .ZN(n36) );
  AOI22_X1 U29 ( .A1(n80), .A2(IN4[10]), .B1(n12), .B2(IN1[9]), .ZN(n35) );
  NAND2_X1 U30 ( .A1(n36), .A2(n35), .ZN(Y[10]) );
  AOI22_X1 U31 ( .A1(n14), .A2(IN4[12]), .B1(n21), .B2(IN1[11]), .ZN(n38) );
  AOI22_X1 U32 ( .A1(n80), .A2(IN4[11]), .B1(n12), .B2(IN1[10]), .ZN(n37) );
  NAND2_X1 U33 ( .A1(n38), .A2(n37), .ZN(Y[11]) );
  AOI22_X1 U34 ( .A1(n14), .A2(IN4[13]), .B1(n21), .B2(IN1[12]), .ZN(n40) );
  AOI22_X1 U35 ( .A1(n80), .A2(IN4[12]), .B1(n12), .B2(IN1[11]), .ZN(n39) );
  NAND2_X1 U36 ( .A1(n40), .A2(n39), .ZN(Y[12]) );
  AOI22_X1 U37 ( .A1(n14), .A2(IN4[14]), .B1(n21), .B2(IN1[13]), .ZN(n42) );
  AOI22_X1 U38 ( .A1(n80), .A2(IN4[13]), .B1(n12), .B2(IN1[12]), .ZN(n41) );
  NAND2_X1 U39 ( .A1(n42), .A2(n41), .ZN(Y[13]) );
  AOI22_X1 U40 ( .A1(n14), .A2(IN4[15]), .B1(n21), .B2(IN1[14]), .ZN(n44) );
  AOI22_X1 U41 ( .A1(n80), .A2(IN4[14]), .B1(n12), .B2(IN1[13]), .ZN(n43) );
  NAND2_X1 U42 ( .A1(n44), .A2(n43), .ZN(Y[14]) );
  AOI22_X1 U43 ( .A1(n14), .A2(IN4[16]), .B1(n21), .B2(IN1[15]), .ZN(n46) );
  AOI22_X1 U44 ( .A1(n80), .A2(IN4[15]), .B1(n12), .B2(IN1[14]), .ZN(n45) );
  NAND2_X1 U45 ( .A1(n46), .A2(n45), .ZN(Y[15]) );
  AOI22_X1 U46 ( .A1(n14), .A2(IN4[17]), .B1(n21), .B2(IN1[16]), .ZN(n48) );
  AOI22_X1 U47 ( .A1(n80), .A2(IN4[16]), .B1(n12), .B2(IN1[15]), .ZN(n47) );
  NAND2_X1 U48 ( .A1(n48), .A2(n47), .ZN(Y[16]) );
  AOI22_X1 U49 ( .A1(n14), .A2(IN4[18]), .B1(n21), .B2(IN1[17]), .ZN(n50) );
  AOI22_X1 U50 ( .A1(n80), .A2(IN4[17]), .B1(n12), .B2(IN1[16]), .ZN(n49) );
  NAND2_X1 U51 ( .A1(n50), .A2(n49), .ZN(Y[17]) );
  AOI22_X1 U52 ( .A1(n14), .A2(IN4[19]), .B1(n21), .B2(IN1[18]), .ZN(n52) );
  AOI22_X1 U53 ( .A1(n80), .A2(IN4[18]), .B1(n12), .B2(IN1[17]), .ZN(n51) );
  NAND2_X1 U54 ( .A1(n52), .A2(n51), .ZN(Y[18]) );
  AOI22_X1 U55 ( .A1(n14), .A2(IN4[20]), .B1(n21), .B2(IN1[19]), .ZN(n54) );
  AOI22_X1 U56 ( .A1(n80), .A2(IN4[19]), .B1(n12), .B2(IN1[18]), .ZN(n53) );
  NAND2_X1 U57 ( .A1(n54), .A2(n53), .ZN(Y[19]) );
  AOI22_X1 U58 ( .A1(n14), .A2(IN4[21]), .B1(n21), .B2(IN1[20]), .ZN(n56) );
  AOI22_X1 U59 ( .A1(n80), .A2(IN4[20]), .B1(n12), .B2(IN1[19]), .ZN(n55) );
  NAND2_X1 U60 ( .A1(n56), .A2(n55), .ZN(Y[20]) );
  AOI22_X1 U61 ( .A1(n14), .A2(IN4[22]), .B1(n77), .B2(IN1[21]), .ZN(n58) );
  AOI22_X1 U62 ( .A1(n80), .A2(IN4[21]), .B1(n12), .B2(IN1[20]), .ZN(n57) );
  NAND2_X1 U63 ( .A1(n58), .A2(n57), .ZN(Y[21]) );
  AOI22_X1 U64 ( .A1(n14), .A2(IN4[23]), .B1(n77), .B2(IN1[22]), .ZN(n60) );
  AOI22_X1 U65 ( .A1(n80), .A2(IN4[22]), .B1(n12), .B2(IN1[21]), .ZN(n59) );
  NAND2_X1 U66 ( .A1(n60), .A2(n59), .ZN(Y[22]) );
  AOI22_X1 U67 ( .A1(n14), .A2(IN4[24]), .B1(n21), .B2(IN1[23]), .ZN(n62) );
  AOI22_X1 U68 ( .A1(n80), .A2(IN4[23]), .B1(n12), .B2(IN1[22]), .ZN(n61) );
  NAND2_X1 U69 ( .A1(n62), .A2(n61), .ZN(Y[23]) );
  AOI22_X1 U70 ( .A1(n14), .A2(IN4[25]), .B1(n21), .B2(IN1[24]), .ZN(n64) );
  AOI22_X1 U71 ( .A1(n80), .A2(IN4[24]), .B1(n12), .B2(IN1[23]), .ZN(n63) );
  NAND2_X1 U72 ( .A1(n64), .A2(n63), .ZN(Y[24]) );
  AOI22_X1 U73 ( .A1(n14), .A2(IN4[26]), .B1(n21), .B2(IN1[25]), .ZN(n66) );
  AOI22_X1 U74 ( .A1(n80), .A2(IN4[25]), .B1(n12), .B2(IN1[24]), .ZN(n65) );
  NAND2_X1 U75 ( .A1(n66), .A2(n65), .ZN(Y[25]) );
  AOI22_X1 U76 ( .A1(n14), .A2(IN4[27]), .B1(n21), .B2(IN1[26]), .ZN(n68) );
  AOI22_X1 U77 ( .A1(n80), .A2(IN4[26]), .B1(n12), .B2(IN1[25]), .ZN(n67) );
  AOI22_X1 U78 ( .A1(n14), .A2(IN4[28]), .B1(n21), .B2(IN1[27]), .ZN(n70) );
  AOI22_X1 U79 ( .A1(n80), .A2(IN4[27]), .B1(n12), .B2(IN1[26]), .ZN(n69) );
  NAND2_X1 U80 ( .A1(n70), .A2(n69), .ZN(Y[27]) );
  AOI22_X1 U81 ( .A1(n14), .A2(IN4[29]), .B1(n21), .B2(IN1[28]), .ZN(n72) );
  AOI22_X1 U82 ( .A1(n80), .A2(IN4[28]), .B1(n12), .B2(IN1[27]), .ZN(n71) );
  NAND2_X1 U83 ( .A1(n72), .A2(n71), .ZN(Y[28]) );
  AOI22_X1 U84 ( .A1(n14), .A2(IN4[30]), .B1(n21), .B2(IN1[29]), .ZN(n74) );
  AOI22_X1 U85 ( .A1(n80), .A2(IN4[29]), .B1(n12), .B2(IN1[28]), .ZN(n73) );
  NAND2_X1 U86 ( .A1(n74), .A2(n73), .ZN(Y[29]) );
  AOI22_X1 U87 ( .A1(n14), .A2(IN4[31]), .B1(n21), .B2(IN1[30]), .ZN(n76) );
  AOI22_X1 U88 ( .A1(n80), .A2(IN4[30]), .B1(n12), .B2(IN1[29]), .ZN(n75) );
  NAND2_X1 U89 ( .A1(n76), .A2(n75), .ZN(Y[30]) );
  AOI22_X1 U90 ( .A1(n14), .A2(IN2[31]), .B1(n21), .B2(IN1[31]), .ZN(n82) );
  AOI22_X1 U91 ( .A1(n80), .A2(IN4[31]), .B1(n12), .B2(IN1[30]), .ZN(n81) );
  NAND2_X1 U92 ( .A1(n82), .A2(n81), .ZN(Y[31]) );
endmodule


module MUX_8to1_N64_13 ( IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, SEL, Y );
  input [63:0] IN0;
  input [63:0] IN1;
  input [63:0] IN2;
  input [63:0] IN3;
  input [63:0] IN4;
  input [63:0] IN5;
  input [63:0] IN6;
  input [63:0] IN7;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n12, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78;

  AND3_X2 U1 ( .A1(n24), .A2(n23), .A3(SEL[2]), .ZN(n76) );
  NAND2_X1 U2 ( .A1(n56), .A2(n55), .ZN(Y[22]) );
  BUF_X1 U3 ( .A(n75), .Z(n21) );
  BUF_X1 U4 ( .A(n73), .Z(n20) );
  BUF_X2 U5 ( .A(n74), .Z(n12) );
  INV_X1 U6 ( .A(SEL[1]), .ZN(n24) );
  NOR3_X1 U7 ( .A1(SEL[2]), .A2(SEL[0]), .A3(n24), .ZN(n74) );
  INV_X1 U8 ( .A(SEL[0]), .ZN(n23) );
  NOR3_X1 U9 ( .A1(SEL[2]), .A2(SEL[1]), .A3(n23), .ZN(n73) );
  OAI21_X1 U10 ( .B1(n12), .B2(n20), .A(IN1[6]), .ZN(n22) );
  INV_X1 U11 ( .A(n22), .ZN(Y[6]) );
  NOR3_X1 U12 ( .A1(SEL[2]), .A2(n24), .A3(n23), .ZN(n75) );
  OAI21_X1 U13 ( .B1(n76), .B2(n21), .A(IN1[6]), .ZN(n26) );
  AOI22_X1 U14 ( .A1(n12), .A2(IN4[8]), .B1(n20), .B2(IN1[7]), .ZN(n25) );
  NAND2_X1 U15 ( .A1(n26), .A2(n25), .ZN(Y[7]) );
  AOI22_X1 U16 ( .A1(n12), .A2(IN4[9]), .B1(n20), .B2(IN1[8]), .ZN(n28) );
  AOI22_X1 U17 ( .A1(IN4[8]), .A2(n76), .B1(n21), .B2(IN1[7]), .ZN(n27) );
  NAND2_X1 U18 ( .A1(n28), .A2(n27), .ZN(Y[8]) );
  AOI22_X1 U19 ( .A1(n12), .A2(IN4[10]), .B1(n20), .B2(IN1[9]), .ZN(n30) );
  AOI22_X1 U20 ( .A1(n76), .A2(IN4[9]), .B1(n21), .B2(IN1[8]), .ZN(n29) );
  NAND2_X1 U21 ( .A1(n30), .A2(n29), .ZN(Y[9]) );
  AOI22_X1 U22 ( .A1(n12), .A2(IN4[11]), .B1(n20), .B2(IN1[10]), .ZN(n32) );
  AOI22_X1 U23 ( .A1(n76), .A2(IN4[10]), .B1(n21), .B2(IN1[9]), .ZN(n31) );
  NAND2_X1 U24 ( .A1(n32), .A2(n31), .ZN(Y[10]) );
  AOI22_X1 U25 ( .A1(n12), .A2(IN4[12]), .B1(n20), .B2(IN1[11]), .ZN(n34) );
  AOI22_X1 U26 ( .A1(n76), .A2(IN4[11]), .B1(n21), .B2(IN1[10]), .ZN(n33) );
  NAND2_X1 U27 ( .A1(n34), .A2(n33), .ZN(Y[11]) );
  AOI22_X1 U28 ( .A1(n12), .A2(IN4[13]), .B1(n20), .B2(IN1[12]), .ZN(n36) );
  AOI22_X1 U29 ( .A1(n76), .A2(IN4[12]), .B1(n21), .B2(IN1[11]), .ZN(n35) );
  NAND2_X1 U30 ( .A1(n36), .A2(n35), .ZN(Y[12]) );
  AOI22_X1 U31 ( .A1(n12), .A2(IN4[14]), .B1(n20), .B2(IN1[13]), .ZN(n38) );
  AOI22_X1 U32 ( .A1(n76), .A2(IN4[13]), .B1(n21), .B2(IN1[12]), .ZN(n37) );
  NAND2_X1 U33 ( .A1(n38), .A2(n37), .ZN(Y[13]) );
  AOI22_X1 U34 ( .A1(n12), .A2(IN4[15]), .B1(n20), .B2(IN1[14]), .ZN(n40) );
  AOI22_X1 U35 ( .A1(n76), .A2(IN4[14]), .B1(n21), .B2(IN1[13]), .ZN(n39) );
  NAND2_X1 U36 ( .A1(n40), .A2(n39), .ZN(Y[14]) );
  AOI22_X1 U37 ( .A1(n12), .A2(IN4[16]), .B1(n20), .B2(IN1[15]), .ZN(n42) );
  AOI22_X1 U38 ( .A1(n76), .A2(IN4[15]), .B1(n21), .B2(IN1[14]), .ZN(n41) );
  NAND2_X1 U39 ( .A1(n42), .A2(n41), .ZN(Y[15]) );
  AOI22_X1 U40 ( .A1(n12), .A2(IN4[17]), .B1(n20), .B2(IN1[16]), .ZN(n44) );
  AOI22_X1 U41 ( .A1(n76), .A2(IN4[16]), .B1(n21), .B2(IN1[15]), .ZN(n43) );
  NAND2_X1 U42 ( .A1(n44), .A2(n43), .ZN(Y[16]) );
  AOI22_X1 U43 ( .A1(n12), .A2(IN4[18]), .B1(n20), .B2(IN1[17]), .ZN(n46) );
  AOI22_X1 U44 ( .A1(n76), .A2(IN4[17]), .B1(n21), .B2(IN1[16]), .ZN(n45) );
  NAND2_X1 U45 ( .A1(n46), .A2(n45), .ZN(Y[17]) );
  AOI22_X1 U46 ( .A1(n12), .A2(IN4[19]), .B1(n20), .B2(IN1[18]), .ZN(n48) );
  AOI22_X1 U47 ( .A1(n76), .A2(IN4[18]), .B1(n21), .B2(IN1[17]), .ZN(n47) );
  NAND2_X1 U48 ( .A1(n48), .A2(n47), .ZN(Y[18]) );
  AOI22_X1 U49 ( .A1(n12), .A2(IN4[20]), .B1(n20), .B2(IN1[19]), .ZN(n50) );
  AOI22_X1 U50 ( .A1(n76), .A2(IN4[19]), .B1(n21), .B2(IN1[18]), .ZN(n49) );
  NAND2_X1 U51 ( .A1(n50), .A2(n49), .ZN(Y[19]) );
  AOI22_X1 U52 ( .A1(n12), .A2(IN4[21]), .B1(n20), .B2(IN1[20]), .ZN(n52) );
  AOI22_X1 U53 ( .A1(n76), .A2(IN4[20]), .B1(n21), .B2(IN1[19]), .ZN(n51) );
  NAND2_X1 U54 ( .A1(n52), .A2(n51), .ZN(Y[20]) );
  AOI22_X1 U55 ( .A1(n12), .A2(IN4[22]), .B1(n20), .B2(IN1[21]), .ZN(n54) );
  AOI22_X1 U56 ( .A1(n76), .A2(IN4[21]), .B1(n21), .B2(IN1[20]), .ZN(n53) );
  NAND2_X1 U57 ( .A1(n54), .A2(n53), .ZN(Y[21]) );
  AOI22_X1 U58 ( .A1(n12), .A2(IN4[23]), .B1(n20), .B2(IN1[22]), .ZN(n56) );
  AOI22_X1 U59 ( .A1(n76), .A2(IN4[22]), .B1(n21), .B2(IN1[21]), .ZN(n55) );
  AOI22_X1 U60 ( .A1(n12), .A2(IN4[24]), .B1(n20), .B2(IN1[23]), .ZN(n58) );
  AOI22_X1 U61 ( .A1(n76), .A2(IN4[23]), .B1(n21), .B2(IN1[22]), .ZN(n57) );
  NAND2_X1 U62 ( .A1(n58), .A2(n57), .ZN(Y[23]) );
  AOI22_X1 U63 ( .A1(n12), .A2(IN4[25]), .B1(n20), .B2(IN1[24]), .ZN(n60) );
  AOI22_X1 U64 ( .A1(n76), .A2(IN4[24]), .B1(n21), .B2(IN1[23]), .ZN(n59) );
  NAND2_X1 U65 ( .A1(n60), .A2(n59), .ZN(Y[24]) );
  AOI22_X1 U66 ( .A1(n12), .A2(IN4[26]), .B1(n20), .B2(IN1[25]), .ZN(n62) );
  AOI22_X1 U67 ( .A1(n76), .A2(IN4[25]), .B1(n21), .B2(IN1[24]), .ZN(n61) );
  NAND2_X1 U68 ( .A1(n62), .A2(n61), .ZN(Y[25]) );
  AOI22_X1 U69 ( .A1(n12), .A2(IN4[27]), .B1(n20), .B2(IN1[26]), .ZN(n64) );
  AOI22_X1 U70 ( .A1(n76), .A2(IN4[26]), .B1(n21), .B2(IN1[25]), .ZN(n63) );
  NAND2_X1 U71 ( .A1(n64), .A2(n63), .ZN(Y[26]) );
  AOI22_X1 U72 ( .A1(n12), .A2(IN4[28]), .B1(n73), .B2(IN1[27]), .ZN(n66) );
  AOI22_X1 U73 ( .A1(n76), .A2(IN4[27]), .B1(n75), .B2(IN1[26]), .ZN(n65) );
  NAND2_X1 U74 ( .A1(n66), .A2(n65), .ZN(Y[27]) );
  AOI22_X1 U75 ( .A1(n12), .A2(IN4[29]), .B1(n20), .B2(IN1[28]), .ZN(n68) );
  AOI22_X1 U76 ( .A1(n76), .A2(IN4[28]), .B1(n21), .B2(IN1[27]), .ZN(n67) );
  NAND2_X1 U77 ( .A1(n68), .A2(n67), .ZN(Y[28]) );
  AOI22_X1 U78 ( .A1(n12), .A2(IN4[30]), .B1(n20), .B2(IN1[29]), .ZN(n70) );
  AOI22_X1 U79 ( .A1(n76), .A2(IN4[29]), .B1(n21), .B2(IN1[28]), .ZN(n69) );
  NAND2_X1 U80 ( .A1(n70), .A2(n69), .ZN(Y[29]) );
  AOI22_X1 U81 ( .A1(n12), .A2(IN4[31]), .B1(n20), .B2(IN1[30]), .ZN(n72) );
  AOI22_X1 U82 ( .A1(n76), .A2(IN4[30]), .B1(n21), .B2(IN1[29]), .ZN(n71) );
  NAND2_X1 U83 ( .A1(n72), .A2(n71), .ZN(Y[30]) );
  AOI22_X1 U84 ( .A1(n12), .A2(IN2[31]), .B1(n20), .B2(IN1[31]), .ZN(n78) );
  AOI22_X1 U85 ( .A1(n76), .A2(IN4[31]), .B1(n21), .B2(IN1[30]), .ZN(n77) );
  NAND2_X1 U86 ( .A1(n78), .A2(n77), .ZN(Y[31]) );
endmodule


module MUX_8to1_N64_12 ( IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, SEL, Y );
  input [63:0] IN0;
  input [63:0] IN1;
  input [63:0] IN2;
  input [63:0] IN3;
  input [63:0] IN4;
  input [63:0] IN5;
  input [63:0] IN6;
  input [63:0] IN7;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74;

  NOR3_X1 U1 ( .A1(SEL[2]), .A2(SEL[0]), .A3(n24), .ZN(n70) );
  BUF_X1 U2 ( .A(n71), .Z(n19) );
  BUF_X1 U3 ( .A(n70), .Z(n21) );
  BUF_X1 U4 ( .A(n69), .Z(n20) );
  AND3_X1 U5 ( .A1(n24), .A2(n23), .A3(SEL[2]), .ZN(n72) );
  NOR3_X1 U6 ( .A1(SEL[2]), .A2(SEL[1]), .A3(n23), .ZN(n69) );
  NAND2_X1 U7 ( .A1(n68), .A2(n67), .ZN(Y[30]) );
  NAND2_X1 U8 ( .A1(n66), .A2(n65), .ZN(Y[29]) );
  INV_X1 U9 ( .A(SEL[1]), .ZN(n24) );
  INV_X1 U10 ( .A(SEL[0]), .ZN(n23) );
  OAI21_X1 U11 ( .B1(n21), .B2(n69), .A(IN1[8]), .ZN(n22) );
  INV_X1 U12 ( .A(n22), .ZN(Y[8]) );
  NOR3_X1 U13 ( .A1(SEL[2]), .A2(n24), .A3(n23), .ZN(n71) );
  OAI21_X1 U14 ( .B1(n72), .B2(n71), .A(IN1[8]), .ZN(n26) );
  AOI22_X1 U15 ( .A1(n21), .A2(IN4[10]), .B1(n20), .B2(IN1[9]), .ZN(n25) );
  NAND2_X1 U16 ( .A1(n26), .A2(n25), .ZN(Y[9]) );
  AOI22_X1 U17 ( .A1(n21), .A2(IN4[11]), .B1(n20), .B2(IN1[10]), .ZN(n28) );
  AOI22_X1 U18 ( .A1(IN4[10]), .A2(n72), .B1(n71), .B2(IN1[9]), .ZN(n27) );
  NAND2_X1 U19 ( .A1(n28), .A2(n27), .ZN(Y[10]) );
  AOI22_X1 U20 ( .A1(n21), .A2(IN4[12]), .B1(n20), .B2(IN1[11]), .ZN(n30) );
  AOI22_X1 U21 ( .A1(n72), .A2(IN4[11]), .B1(n19), .B2(IN1[10]), .ZN(n29) );
  NAND2_X1 U22 ( .A1(n30), .A2(n29), .ZN(Y[11]) );
  AOI22_X1 U23 ( .A1(n21), .A2(IN4[13]), .B1(n20), .B2(IN1[12]), .ZN(n32) );
  AOI22_X1 U24 ( .A1(n72), .A2(IN4[12]), .B1(n71), .B2(IN1[11]), .ZN(n31) );
  NAND2_X1 U25 ( .A1(n32), .A2(n31), .ZN(Y[12]) );
  AOI22_X1 U26 ( .A1(n21), .A2(IN4[14]), .B1(n20), .B2(IN1[13]), .ZN(n34) );
  AOI22_X1 U27 ( .A1(n72), .A2(IN4[13]), .B1(n19), .B2(IN1[12]), .ZN(n33) );
  NAND2_X1 U28 ( .A1(n34), .A2(n33), .ZN(Y[13]) );
  AOI22_X1 U29 ( .A1(n21), .A2(IN4[15]), .B1(n20), .B2(IN1[14]), .ZN(n36) );
  AOI22_X1 U30 ( .A1(n72), .A2(IN4[14]), .B1(n71), .B2(IN1[13]), .ZN(n35) );
  NAND2_X1 U31 ( .A1(n36), .A2(n35), .ZN(Y[14]) );
  AOI22_X1 U32 ( .A1(n21), .A2(IN4[16]), .B1(n20), .B2(IN1[15]), .ZN(n38) );
  AOI22_X1 U33 ( .A1(n72), .A2(IN4[15]), .B1(n19), .B2(IN1[14]), .ZN(n37) );
  NAND2_X1 U34 ( .A1(n38), .A2(n37), .ZN(Y[15]) );
  AOI22_X1 U35 ( .A1(n21), .A2(IN4[17]), .B1(n20), .B2(IN1[16]), .ZN(n40) );
  AOI22_X1 U36 ( .A1(n72), .A2(IN4[16]), .B1(n19), .B2(IN1[15]), .ZN(n39) );
  NAND2_X1 U37 ( .A1(n40), .A2(n39), .ZN(Y[16]) );
  AOI22_X1 U38 ( .A1(n21), .A2(IN4[18]), .B1(n20), .B2(IN1[17]), .ZN(n42) );
  AOI22_X1 U39 ( .A1(n72), .A2(IN4[17]), .B1(n71), .B2(IN1[16]), .ZN(n41) );
  NAND2_X1 U40 ( .A1(n42), .A2(n41), .ZN(Y[17]) );
  AOI22_X1 U41 ( .A1(n21), .A2(IN4[19]), .B1(n20), .B2(IN1[18]), .ZN(n44) );
  AOI22_X1 U42 ( .A1(n72), .A2(IN4[18]), .B1(n19), .B2(IN1[17]), .ZN(n43) );
  NAND2_X1 U43 ( .A1(n44), .A2(n43), .ZN(Y[18]) );
  AOI22_X1 U44 ( .A1(n21), .A2(IN4[20]), .B1(n20), .B2(IN1[19]), .ZN(n46) );
  AOI22_X1 U45 ( .A1(n72), .A2(IN4[19]), .B1(n71), .B2(IN1[18]), .ZN(n45) );
  NAND2_X1 U46 ( .A1(n46), .A2(n45), .ZN(Y[19]) );
  AOI22_X1 U47 ( .A1(n21), .A2(IN4[21]), .B1(n20), .B2(IN1[20]), .ZN(n48) );
  AOI22_X1 U48 ( .A1(n72), .A2(IN4[20]), .B1(n19), .B2(IN1[19]), .ZN(n47) );
  NAND2_X1 U49 ( .A1(n48), .A2(n47), .ZN(Y[20]) );
  AOI22_X1 U50 ( .A1(n21), .A2(IN4[22]), .B1(n69), .B2(IN1[21]), .ZN(n50) );
  AOI22_X1 U51 ( .A1(n72), .A2(IN4[21]), .B1(n19), .B2(IN1[20]), .ZN(n49) );
  NAND2_X1 U52 ( .A1(n50), .A2(n49), .ZN(Y[21]) );
  AOI22_X1 U53 ( .A1(n21), .A2(IN4[23]), .B1(n69), .B2(IN1[22]), .ZN(n52) );
  AOI22_X1 U54 ( .A1(n72), .A2(IN4[22]), .B1(n19), .B2(IN1[21]), .ZN(n51) );
  NAND2_X1 U55 ( .A1(n52), .A2(n51), .ZN(Y[22]) );
  AOI22_X1 U56 ( .A1(n21), .A2(IN4[24]), .B1(n20), .B2(IN1[23]), .ZN(n54) );
  AOI22_X1 U57 ( .A1(n72), .A2(IN4[23]), .B1(n19), .B2(IN1[22]), .ZN(n53) );
  NAND2_X1 U58 ( .A1(n54), .A2(n53), .ZN(Y[23]) );
  AOI22_X1 U59 ( .A1(n70), .A2(IN4[25]), .B1(n69), .B2(IN1[24]), .ZN(n56) );
  AOI22_X1 U60 ( .A1(n72), .A2(IN4[24]), .B1(n19), .B2(IN1[23]), .ZN(n55) );
  NAND2_X1 U61 ( .A1(n56), .A2(n55), .ZN(Y[24]) );
  AOI22_X1 U62 ( .A1(n21), .A2(IN4[26]), .B1(n69), .B2(IN1[25]), .ZN(n58) );
  AOI22_X1 U63 ( .A1(n72), .A2(IN4[25]), .B1(n19), .B2(IN1[24]), .ZN(n57) );
  NAND2_X1 U64 ( .A1(n58), .A2(n57), .ZN(Y[25]) );
  AOI22_X1 U65 ( .A1(n70), .A2(IN4[27]), .B1(n69), .B2(IN1[26]), .ZN(n60) );
  AOI22_X1 U66 ( .A1(n72), .A2(IN4[26]), .B1(n19), .B2(IN1[25]), .ZN(n59) );
  NAND2_X1 U67 ( .A1(n60), .A2(n59), .ZN(Y[26]) );
  AOI22_X1 U68 ( .A1(n70), .A2(IN4[28]), .B1(n20), .B2(IN1[27]), .ZN(n62) );
  AOI22_X1 U69 ( .A1(n72), .A2(IN4[27]), .B1(n19), .B2(IN1[26]), .ZN(n61) );
  NAND2_X1 U70 ( .A1(n62), .A2(n61), .ZN(Y[27]) );
  AOI22_X1 U71 ( .A1(n70), .A2(IN4[29]), .B1(n20), .B2(IN1[28]), .ZN(n64) );
  AOI22_X1 U72 ( .A1(n72), .A2(IN4[28]), .B1(n19), .B2(IN1[27]), .ZN(n63) );
  NAND2_X1 U73 ( .A1(n64), .A2(n63), .ZN(Y[28]) );
  AOI22_X1 U74 ( .A1(n70), .A2(IN4[30]), .B1(n20), .B2(IN1[29]), .ZN(n66) );
  AOI22_X1 U75 ( .A1(n72), .A2(IN4[29]), .B1(n19), .B2(IN1[28]), .ZN(n65) );
  AOI22_X1 U76 ( .A1(n70), .A2(IN4[31]), .B1(n20), .B2(IN1[30]), .ZN(n68) );
  AOI22_X1 U77 ( .A1(n72), .A2(IN4[30]), .B1(n19), .B2(IN1[29]), .ZN(n67) );
  AOI22_X1 U78 ( .A1(n21), .A2(IN2[31]), .B1(n20), .B2(IN1[31]), .ZN(n74) );
  AOI22_X1 U79 ( .A1(n72), .A2(IN4[31]), .B1(n19), .B2(IN1[30]), .ZN(n73) );
  NAND2_X1 U80 ( .A1(n74), .A2(n73), .ZN(Y[31]) );
endmodule


module MUX_8to1_N64_11 ( IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, SEL, Y );
  input [63:0] IN0;
  input [63:0] IN1;
  input [63:0] IN2;
  input [63:0] IN3;
  input [63:0] IN4;
  input [63:0] IN5;
  input [63:0] IN6;
  input [63:0] IN7;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n4, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70;

  CLKBUF_X3 U1 ( .A(n66), .Z(n19) );
  CLKBUF_X3 U2 ( .A(n67), .Z(n21) );
  BUF_X2 U3 ( .A(n65), .Z(n4) );
  CLKBUF_X3 U4 ( .A(n66), .Z(n18) );
  CLKBUF_X3 U5 ( .A(n67), .Z(n20) );
  AND3_X2 U6 ( .A1(n24), .A2(n23), .A3(SEL[2]), .ZN(n68) );
  INV_X1 U7 ( .A(SEL[1]), .ZN(n24) );
  NOR3_X1 U8 ( .A1(SEL[2]), .A2(SEL[0]), .A3(n24), .ZN(n66) );
  INV_X1 U9 ( .A(SEL[0]), .ZN(n23) );
  NOR3_X1 U10 ( .A1(SEL[2]), .A2(n23), .A3(SEL[1]), .ZN(n65) );
  OAI21_X1 U11 ( .B1(n19), .B2(n4), .A(IN1[10]), .ZN(n22) );
  INV_X1 U12 ( .A(n22), .ZN(Y[10]) );
  NOR3_X1 U13 ( .A1(SEL[2]), .A2(n24), .A3(n23), .ZN(n67) );
  OAI21_X1 U14 ( .B1(n68), .B2(n21), .A(IN1[10]), .ZN(n26) );
  AOI22_X1 U15 ( .A1(n18), .A2(IN4[12]), .B1(n4), .B2(IN1[11]), .ZN(n25) );
  NAND2_X1 U16 ( .A1(n26), .A2(n25), .ZN(Y[11]) );
  AOI22_X1 U17 ( .A1(n19), .A2(IN4[13]), .B1(n4), .B2(IN1[12]), .ZN(n28) );
  AOI22_X1 U18 ( .A1(IN4[12]), .A2(n68), .B1(n20), .B2(IN1[11]), .ZN(n27) );
  NAND2_X1 U19 ( .A1(n28), .A2(n27), .ZN(Y[12]) );
  AOI22_X1 U20 ( .A1(n19), .A2(IN4[14]), .B1(n4), .B2(IN1[13]), .ZN(n30) );
  AOI22_X1 U21 ( .A1(n68), .A2(IN4[13]), .B1(n20), .B2(IN1[12]), .ZN(n29) );
  NAND2_X1 U22 ( .A1(n30), .A2(n29), .ZN(Y[13]) );
  AOI22_X1 U23 ( .A1(n18), .A2(IN4[15]), .B1(n4), .B2(IN1[14]), .ZN(n32) );
  AOI22_X1 U24 ( .A1(n68), .A2(IN4[14]), .B1(n21), .B2(IN1[13]), .ZN(n31) );
  NAND2_X1 U25 ( .A1(n32), .A2(n31), .ZN(Y[14]) );
  AOI22_X1 U26 ( .A1(n18), .A2(IN4[16]), .B1(n4), .B2(IN1[15]), .ZN(n34) );
  AOI22_X1 U27 ( .A1(n68), .A2(IN4[15]), .B1(n21), .B2(IN1[14]), .ZN(n33) );
  NAND2_X1 U28 ( .A1(n34), .A2(n33), .ZN(Y[15]) );
  AOI22_X1 U29 ( .A1(n19), .A2(IN4[17]), .B1(n4), .B2(IN1[16]), .ZN(n36) );
  AOI22_X1 U30 ( .A1(n68), .A2(IN4[16]), .B1(n21), .B2(IN1[15]), .ZN(n35) );
  NAND2_X1 U31 ( .A1(n36), .A2(n35), .ZN(Y[16]) );
  AOI22_X1 U32 ( .A1(n19), .A2(IN4[18]), .B1(n4), .B2(IN1[17]), .ZN(n38) );
  AOI22_X1 U33 ( .A1(n68), .A2(IN4[17]), .B1(n20), .B2(IN1[16]), .ZN(n37) );
  NAND2_X1 U34 ( .A1(n38), .A2(n37), .ZN(Y[17]) );
  AOI22_X1 U35 ( .A1(n18), .A2(IN4[19]), .B1(n4), .B2(IN1[18]), .ZN(n40) );
  AOI22_X1 U36 ( .A1(n68), .A2(IN4[18]), .B1(n20), .B2(IN1[17]), .ZN(n39) );
  NAND2_X1 U37 ( .A1(n40), .A2(n39), .ZN(Y[18]) );
  AOI22_X1 U38 ( .A1(n18), .A2(IN4[20]), .B1(n4), .B2(IN1[19]), .ZN(n42) );
  AOI22_X1 U39 ( .A1(n68), .A2(IN4[19]), .B1(n21), .B2(IN1[18]), .ZN(n41) );
  NAND2_X1 U40 ( .A1(n42), .A2(n41), .ZN(Y[19]) );
  AOI22_X1 U41 ( .A1(IN4[21]), .A2(n19), .B1(n4), .B2(IN1[20]), .ZN(n44) );
  AOI22_X1 U42 ( .A1(n68), .A2(IN4[20]), .B1(n20), .B2(IN1[19]), .ZN(n43) );
  NAND2_X1 U43 ( .A1(n44), .A2(n43), .ZN(Y[20]) );
  AOI22_X1 U44 ( .A1(n19), .A2(IN4[22]), .B1(n4), .B2(IN1[21]), .ZN(n46) );
  AOI22_X1 U45 ( .A1(n68), .A2(IN4[21]), .B1(n20), .B2(IN1[20]), .ZN(n45) );
  NAND2_X1 U46 ( .A1(n46), .A2(n45), .ZN(Y[21]) );
  AOI22_X1 U47 ( .A1(n18), .A2(IN4[23]), .B1(n4), .B2(IN1[22]), .ZN(n48) );
  AOI22_X1 U48 ( .A1(n68), .A2(IN4[22]), .B1(n20), .B2(IN1[21]), .ZN(n47) );
  NAND2_X1 U49 ( .A1(n48), .A2(n47), .ZN(Y[22]) );
  AOI22_X1 U50 ( .A1(n18), .A2(IN4[24]), .B1(n4), .B2(IN1[23]), .ZN(n50) );
  AOI22_X1 U51 ( .A1(n68), .A2(IN4[23]), .B1(n21), .B2(IN1[22]), .ZN(n49) );
  NAND2_X1 U52 ( .A1(n50), .A2(n49), .ZN(Y[23]) );
  AOI22_X1 U53 ( .A1(n19), .A2(IN4[25]), .B1(n4), .B2(IN1[24]), .ZN(n52) );
  AOI22_X1 U54 ( .A1(n68), .A2(IN4[24]), .B1(n21), .B2(IN1[23]), .ZN(n51) );
  NAND2_X1 U55 ( .A1(n52), .A2(n51), .ZN(Y[24]) );
  AOI22_X1 U56 ( .A1(n19), .A2(IN4[26]), .B1(n4), .B2(IN1[25]), .ZN(n54) );
  AOI22_X1 U57 ( .A1(n68), .A2(IN4[25]), .B1(n21), .B2(IN1[24]), .ZN(n53) );
  NAND2_X1 U58 ( .A1(n54), .A2(n53), .ZN(Y[25]) );
  AOI22_X1 U59 ( .A1(n18), .A2(IN4[27]), .B1(n4), .B2(IN1[26]), .ZN(n56) );
  AOI22_X1 U60 ( .A1(n68), .A2(IN4[26]), .B1(n20), .B2(IN1[25]), .ZN(n55) );
  NAND2_X1 U61 ( .A1(n56), .A2(n55), .ZN(Y[26]) );
  AOI22_X1 U62 ( .A1(n18), .A2(IN4[28]), .B1(n4), .B2(IN1[27]), .ZN(n58) );
  AOI22_X1 U63 ( .A1(n68), .A2(IN4[27]), .B1(n20), .B2(IN1[26]), .ZN(n57) );
  NAND2_X1 U64 ( .A1(n58), .A2(n57), .ZN(Y[27]) );
  AOI22_X1 U65 ( .A1(n19), .A2(IN4[29]), .B1(n4), .B2(IN1[28]), .ZN(n60) );
  AOI22_X1 U66 ( .A1(n68), .A2(IN4[28]), .B1(n21), .B2(IN1[27]), .ZN(n59) );
  NAND2_X1 U67 ( .A1(n60), .A2(n59), .ZN(Y[28]) );
  AOI22_X1 U68 ( .A1(n19), .A2(IN4[30]), .B1(n4), .B2(IN1[29]), .ZN(n62) );
  AOI22_X1 U69 ( .A1(n68), .A2(IN4[29]), .B1(n20), .B2(IN1[28]), .ZN(n61) );
  NAND2_X1 U70 ( .A1(n62), .A2(n61), .ZN(Y[29]) );
  AOI22_X1 U71 ( .A1(n18), .A2(IN4[31]), .B1(n4), .B2(IN1[30]), .ZN(n64) );
  AOI22_X1 U72 ( .A1(n68), .A2(IN4[30]), .B1(n21), .B2(IN1[29]), .ZN(n63) );
  NAND2_X1 U73 ( .A1(n64), .A2(n63), .ZN(Y[30]) );
  AOI22_X1 U74 ( .A1(n18), .A2(IN2[31]), .B1(n4), .B2(IN1[31]), .ZN(n70) );
  AOI22_X1 U75 ( .A1(n68), .A2(IN4[31]), .B1(n20), .B2(IN1[30]), .ZN(n69) );
  NAND2_X1 U76 ( .A1(n70), .A2(n69), .ZN(Y[31]) );
endmodule


module MUX_8to1_N64_10 ( IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, SEL, Y );
  input [63:0] IN0;
  input [63:0] IN1;
  input [63:0] IN2;
  input [63:0] IN3;
  input [63:0] IN4;
  input [63:0] IN5;
  input [63:0] IN6;
  input [63:0] IN7;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62;

  BUF_X1 U1 ( .A(n58), .Z(n16) );
  BUF_X1 U2 ( .A(n57), .Z(n17) );
  AND3_X1 U3 ( .A1(n20), .A2(n19), .A3(SEL[2]), .ZN(n60) );
  NOR3_X4 U4 ( .A1(SEL[2]), .A2(n20), .A3(n19), .ZN(n59) );
  INV_X1 U5 ( .A(SEL[1]), .ZN(n20) );
  NOR3_X1 U6 ( .A1(SEL[2]), .A2(SEL[1]), .A3(n19), .ZN(n57) );
  NOR3_X1 U7 ( .A1(SEL[2]), .A2(SEL[0]), .A3(n20), .ZN(n58) );
  INV_X1 U8 ( .A(SEL[0]), .ZN(n19) );
  OAI21_X1 U9 ( .B1(n16), .B2(n17), .A(IN1[12]), .ZN(n18) );
  INV_X1 U10 ( .A(n18), .ZN(Y[12]) );
  OAI21_X1 U11 ( .B1(n60), .B2(n59), .A(IN1[12]), .ZN(n22) );
  AOI22_X1 U12 ( .A1(n16), .A2(IN4[14]), .B1(n57), .B2(IN1[13]), .ZN(n21) );
  NAND2_X1 U13 ( .A1(n22), .A2(n21), .ZN(Y[13]) );
  AOI22_X1 U14 ( .A1(n16), .A2(IN4[15]), .B1(n57), .B2(IN1[14]), .ZN(n24) );
  AOI22_X1 U15 ( .A1(n60), .A2(IN4[14]), .B1(n59), .B2(IN1[13]), .ZN(n23) );
  NAND2_X1 U16 ( .A1(n24), .A2(n23), .ZN(Y[14]) );
  AOI22_X1 U17 ( .A1(n16), .A2(IN4[16]), .B1(n17), .B2(IN1[15]), .ZN(n26) );
  AOI22_X1 U18 ( .A1(n60), .A2(IN4[15]), .B1(n59), .B2(IN1[14]), .ZN(n25) );
  NAND2_X1 U19 ( .A1(n26), .A2(n25), .ZN(Y[15]) );
  AOI22_X1 U20 ( .A1(n16), .A2(IN4[17]), .B1(n17), .B2(IN1[16]), .ZN(n28) );
  AOI22_X1 U21 ( .A1(n60), .A2(IN4[16]), .B1(n59), .B2(IN1[15]), .ZN(n27) );
  NAND2_X1 U22 ( .A1(n28), .A2(n27), .ZN(Y[16]) );
  AOI22_X1 U23 ( .A1(n16), .A2(IN4[18]), .B1(n57), .B2(IN1[17]), .ZN(n30) );
  AOI22_X1 U24 ( .A1(n60), .A2(IN4[17]), .B1(n59), .B2(IN1[16]), .ZN(n29) );
  NAND2_X1 U25 ( .A1(n30), .A2(n29), .ZN(Y[17]) );
  AOI22_X1 U26 ( .A1(n16), .A2(IN4[19]), .B1(n57), .B2(IN1[18]), .ZN(n32) );
  AOI22_X1 U27 ( .A1(n60), .A2(IN4[18]), .B1(n59), .B2(IN1[17]), .ZN(n31) );
  NAND2_X1 U28 ( .A1(n32), .A2(n31), .ZN(Y[18]) );
  AOI22_X1 U29 ( .A1(n16), .A2(IN4[20]), .B1(n17), .B2(IN1[19]), .ZN(n34) );
  AOI22_X1 U30 ( .A1(n60), .A2(IN4[19]), .B1(n59), .B2(IN1[18]), .ZN(n33) );
  NAND2_X1 U31 ( .A1(n34), .A2(n33), .ZN(Y[19]) );
  AOI22_X1 U32 ( .A1(n16), .A2(IN4[21]), .B1(n17), .B2(IN1[20]), .ZN(n36) );
  AOI22_X1 U33 ( .A1(n60), .A2(IN4[20]), .B1(n59), .B2(IN1[19]), .ZN(n35) );
  NAND2_X1 U34 ( .A1(n36), .A2(n35), .ZN(Y[20]) );
  AOI22_X1 U35 ( .A1(n16), .A2(IN4[22]), .B1(n17), .B2(IN1[21]), .ZN(n38) );
  AOI22_X1 U36 ( .A1(n60), .A2(IN4[21]), .B1(n59), .B2(IN1[20]), .ZN(n37) );
  NAND2_X1 U37 ( .A1(n38), .A2(n37), .ZN(Y[21]) );
  AOI22_X1 U38 ( .A1(n16), .A2(IN4[23]), .B1(n17), .B2(IN1[22]), .ZN(n40) );
  AOI22_X1 U39 ( .A1(n60), .A2(IN4[22]), .B1(n59), .B2(IN1[21]), .ZN(n39) );
  NAND2_X1 U40 ( .A1(n40), .A2(n39), .ZN(Y[22]) );
  AOI22_X1 U41 ( .A1(n16), .A2(IN4[24]), .B1(n17), .B2(IN1[23]), .ZN(n42) );
  AOI22_X1 U42 ( .A1(n60), .A2(IN4[23]), .B1(n59), .B2(IN1[22]), .ZN(n41) );
  NAND2_X1 U43 ( .A1(n42), .A2(n41), .ZN(Y[23]) );
  AOI22_X1 U44 ( .A1(n58), .A2(IN4[25]), .B1(n17), .B2(IN1[24]), .ZN(n44) );
  AOI22_X1 U45 ( .A1(n60), .A2(IN4[24]), .B1(n59), .B2(IN1[23]), .ZN(n43) );
  NAND2_X1 U46 ( .A1(n44), .A2(n43), .ZN(Y[24]) );
  AOI22_X1 U47 ( .A1(n16), .A2(IN4[26]), .B1(n17), .B2(IN1[25]), .ZN(n46) );
  AOI22_X1 U48 ( .A1(n60), .A2(IN4[25]), .B1(n59), .B2(IN1[24]), .ZN(n45) );
  NAND2_X1 U49 ( .A1(n46), .A2(n45), .ZN(Y[25]) );
  AOI22_X1 U50 ( .A1(n16), .A2(IN4[27]), .B1(n17), .B2(IN1[26]), .ZN(n48) );
  AOI22_X1 U51 ( .A1(n60), .A2(IN4[26]), .B1(n59), .B2(IN1[25]), .ZN(n47) );
  NAND2_X1 U52 ( .A1(n48), .A2(n47), .ZN(Y[26]) );
  AOI22_X1 U53 ( .A1(n58), .A2(IN4[28]), .B1(n57), .B2(IN1[27]), .ZN(n50) );
  AOI22_X1 U54 ( .A1(n60), .A2(IN4[27]), .B1(n59), .B2(IN1[26]), .ZN(n49) );
  NAND2_X1 U55 ( .A1(n50), .A2(n49), .ZN(Y[27]) );
  AOI22_X1 U56 ( .A1(n58), .A2(IN4[29]), .B1(n57), .B2(IN1[28]), .ZN(n52) );
  AOI22_X1 U57 ( .A1(n60), .A2(IN4[28]), .B1(n59), .B2(IN1[27]), .ZN(n51) );
  NAND2_X1 U58 ( .A1(n52), .A2(n51), .ZN(Y[28]) );
  AOI22_X1 U59 ( .A1(n16), .A2(IN4[30]), .B1(n17), .B2(IN1[29]), .ZN(n54) );
  AOI22_X1 U60 ( .A1(n60), .A2(IN4[29]), .B1(n59), .B2(IN1[28]), .ZN(n53) );
  NAND2_X1 U61 ( .A1(n54), .A2(n53), .ZN(Y[29]) );
  AOI22_X1 U62 ( .A1(n16), .A2(IN4[31]), .B1(n17), .B2(IN1[30]), .ZN(n56) );
  AOI22_X1 U63 ( .A1(n60), .A2(IN4[30]), .B1(n59), .B2(IN1[29]), .ZN(n55) );
  NAND2_X1 U64 ( .A1(n56), .A2(n55), .ZN(Y[30]) );
  AOI22_X1 U65 ( .A1(n58), .A2(IN2[31]), .B1(n17), .B2(IN1[31]), .ZN(n62) );
  AOI22_X1 U66 ( .A1(n60), .A2(IN4[31]), .B1(n59), .B2(IN1[30]), .ZN(n61) );
  NAND2_X1 U67 ( .A1(n62), .A2(n61), .ZN(Y[31]) );
endmodule


module MUX_8to1_N64_9 ( IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, SEL, Y );
  input [63:0] IN0;
  input [63:0] IN1;
  input [63:0] IN2;
  input [63:0] IN3;
  input [63:0] IN4;
  input [63:0] IN5;
  input [63:0] IN6;
  input [63:0] IN7;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54;

  INV_X1 U1 ( .A(n51), .ZN(n13) );
  INV_X1 U2 ( .A(n14), .ZN(Y[14]) );
  OR3_X1 U3 ( .A1(SEL[2]), .A2(n16), .A3(n15), .ZN(n51) );
  AND3_X1 U4 ( .A1(n16), .A2(n15), .A3(SEL[2]), .ZN(n52) );
  NOR3_X4 U5 ( .A1(SEL[2]), .A2(SEL[1]), .A3(n15), .ZN(n49) );
  NOR3_X4 U6 ( .A1(SEL[2]), .A2(SEL[0]), .A3(n16), .ZN(n50) );
  INV_X1 U7 ( .A(SEL[1]), .ZN(n16) );
  INV_X1 U8 ( .A(SEL[0]), .ZN(n15) );
  OAI21_X1 U9 ( .B1(n50), .B2(n49), .A(IN1[14]), .ZN(n14) );
  OAI21_X1 U10 ( .B1(n52), .B2(n13), .A(IN1[14]), .ZN(n18) );
  AOI22_X1 U11 ( .A1(n50), .A2(IN4[16]), .B1(n49), .B2(IN1[15]), .ZN(n17) );
  NAND2_X1 U12 ( .A1(n18), .A2(n17), .ZN(Y[15]) );
  AOI22_X1 U13 ( .A1(n50), .A2(IN4[17]), .B1(n49), .B2(IN1[16]), .ZN(n20) );
  AOI22_X1 U14 ( .A1(n52), .A2(IN4[16]), .B1(n13), .B2(IN1[15]), .ZN(n19) );
  NAND2_X1 U15 ( .A1(n20), .A2(n19), .ZN(Y[16]) );
  AOI22_X1 U16 ( .A1(n50), .A2(IN4[18]), .B1(n49), .B2(IN1[17]), .ZN(n22) );
  AOI22_X1 U17 ( .A1(n52), .A2(IN4[17]), .B1(n13), .B2(IN1[16]), .ZN(n21) );
  NAND2_X1 U18 ( .A1(n22), .A2(n21), .ZN(Y[17]) );
  AOI22_X1 U19 ( .A1(n50), .A2(IN4[19]), .B1(n49), .B2(IN1[18]), .ZN(n24) );
  AOI22_X1 U20 ( .A1(n52), .A2(IN4[18]), .B1(n13), .B2(IN1[17]), .ZN(n23) );
  NAND2_X1 U21 ( .A1(n24), .A2(n23), .ZN(Y[18]) );
  AOI22_X1 U22 ( .A1(n50), .A2(IN4[20]), .B1(n49), .B2(IN1[19]), .ZN(n26) );
  AOI22_X1 U23 ( .A1(n52), .A2(IN4[19]), .B1(n13), .B2(IN1[18]), .ZN(n25) );
  NAND2_X1 U24 ( .A1(n26), .A2(n25), .ZN(Y[19]) );
  AOI22_X1 U25 ( .A1(n50), .A2(IN4[21]), .B1(n49), .B2(IN1[20]), .ZN(n28) );
  AOI22_X1 U26 ( .A1(n52), .A2(IN4[20]), .B1(n13), .B2(IN1[19]), .ZN(n27) );
  NAND2_X1 U27 ( .A1(n28), .A2(n27), .ZN(Y[20]) );
  AOI22_X1 U28 ( .A1(n50), .A2(IN4[22]), .B1(n49), .B2(IN1[21]), .ZN(n30) );
  AOI22_X1 U29 ( .A1(n52), .A2(IN4[21]), .B1(n13), .B2(IN1[20]), .ZN(n29) );
  NAND2_X1 U30 ( .A1(n30), .A2(n29), .ZN(Y[21]) );
  AOI22_X1 U31 ( .A1(n50), .A2(IN4[23]), .B1(n49), .B2(IN1[22]), .ZN(n32) );
  AOI22_X1 U32 ( .A1(n52), .A2(IN4[22]), .B1(n13), .B2(IN1[21]), .ZN(n31) );
  NAND2_X1 U33 ( .A1(n32), .A2(n31), .ZN(Y[22]) );
  AOI22_X1 U34 ( .A1(n50), .A2(IN4[24]), .B1(n49), .B2(IN1[23]), .ZN(n34) );
  AOI22_X1 U35 ( .A1(n52), .A2(IN4[23]), .B1(n13), .B2(IN1[22]), .ZN(n33) );
  NAND2_X1 U36 ( .A1(n34), .A2(n33), .ZN(Y[23]) );
  AOI22_X1 U37 ( .A1(n50), .A2(IN4[25]), .B1(n49), .B2(IN1[24]), .ZN(n36) );
  AOI22_X1 U38 ( .A1(n52), .A2(IN4[24]), .B1(n13), .B2(IN1[23]), .ZN(n35) );
  NAND2_X1 U39 ( .A1(n36), .A2(n35), .ZN(Y[24]) );
  AOI22_X1 U40 ( .A1(n50), .A2(IN4[26]), .B1(n49), .B2(IN1[25]), .ZN(n38) );
  AOI22_X1 U41 ( .A1(n52), .A2(IN4[25]), .B1(n13), .B2(IN1[24]), .ZN(n37) );
  NAND2_X1 U42 ( .A1(n38), .A2(n37), .ZN(Y[25]) );
  AOI22_X1 U43 ( .A1(n50), .A2(IN4[27]), .B1(n49), .B2(IN1[26]), .ZN(n40) );
  AOI22_X1 U44 ( .A1(n52), .A2(IN4[26]), .B1(n13), .B2(IN1[25]), .ZN(n39) );
  NAND2_X1 U45 ( .A1(n40), .A2(n39), .ZN(Y[26]) );
  AOI22_X1 U46 ( .A1(n50), .A2(IN4[28]), .B1(n49), .B2(IN1[27]), .ZN(n42) );
  AOI22_X1 U47 ( .A1(n52), .A2(IN4[27]), .B1(n13), .B2(IN1[26]), .ZN(n41) );
  NAND2_X1 U48 ( .A1(n42), .A2(n41), .ZN(Y[27]) );
  AOI22_X1 U49 ( .A1(n50), .A2(IN4[29]), .B1(n49), .B2(IN1[28]), .ZN(n44) );
  AOI22_X1 U50 ( .A1(n52), .A2(IN4[28]), .B1(n13), .B2(IN1[27]), .ZN(n43) );
  NAND2_X1 U51 ( .A1(n44), .A2(n43), .ZN(Y[28]) );
  AOI22_X1 U52 ( .A1(n50), .A2(IN4[30]), .B1(n49), .B2(IN1[29]), .ZN(n46) );
  AOI22_X1 U53 ( .A1(n52), .A2(IN4[29]), .B1(n13), .B2(IN1[28]), .ZN(n45) );
  NAND2_X1 U54 ( .A1(n46), .A2(n45), .ZN(Y[29]) );
  AOI22_X1 U55 ( .A1(n50), .A2(IN4[31]), .B1(n49), .B2(IN1[30]), .ZN(n48) );
  AOI22_X1 U56 ( .A1(n52), .A2(IN4[30]), .B1(n13), .B2(IN1[29]), .ZN(n47) );
  NAND2_X1 U57 ( .A1(n48), .A2(n47), .ZN(Y[30]) );
  AOI22_X1 U58 ( .A1(n50), .A2(IN2[31]), .B1(n49), .B2(IN1[31]), .ZN(n54) );
  AOI22_X1 U59 ( .A1(n52), .A2(IN4[31]), .B1(n13), .B2(IN1[30]), .ZN(n53) );
  NAND2_X1 U60 ( .A1(n54), .A2(n53), .ZN(Y[31]) );
endmodule


module MUX_8to1_N64_8 ( IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, SEL, Y );
  input [63:0] IN0;
  input [63:0] IN1;
  input [63:0] IN2;
  input [63:0] IN3;
  input [63:0] IN4;
  input [63:0] IN5;
  input [63:0] IN6;
  input [63:0] IN7;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50;

  INV_X1 U1 ( .A(n14), .ZN(Y[16]) );
  AND3_X1 U2 ( .A1(n16), .A2(n15), .A3(SEL[2]), .ZN(n48) );
  OR3_X1 U3 ( .A1(SEL[2]), .A2(n16), .A3(n15), .ZN(n47) );
  OR3_X1 U4 ( .A1(SEL[2]), .A2(SEL[1]), .A3(n15), .ZN(n45) );
  INV_X1 U5 ( .A(n47), .ZN(n12) );
  INV_X1 U6 ( .A(n45), .ZN(n13) );
  NOR3_X4 U7 ( .A1(SEL[2]), .A2(SEL[0]), .A3(n16), .ZN(n46) );
  INV_X1 U8 ( .A(SEL[1]), .ZN(n16) );
  INV_X1 U9 ( .A(SEL[0]), .ZN(n15) );
  OAI21_X1 U10 ( .B1(n46), .B2(n13), .A(IN1[16]), .ZN(n14) );
  OAI21_X1 U11 ( .B1(n48), .B2(n12), .A(IN1[16]), .ZN(n18) );
  AOI22_X1 U12 ( .A1(n46), .A2(IN4[18]), .B1(n13), .B2(IN1[17]), .ZN(n17) );
  NAND2_X1 U13 ( .A1(n18), .A2(n17), .ZN(Y[17]) );
  AOI22_X1 U14 ( .A1(n46), .A2(IN4[19]), .B1(n13), .B2(IN1[18]), .ZN(n20) );
  AOI22_X1 U15 ( .A1(n48), .A2(IN4[18]), .B1(n12), .B2(IN1[17]), .ZN(n19) );
  NAND2_X1 U16 ( .A1(n20), .A2(n19), .ZN(Y[18]) );
  AOI22_X1 U17 ( .A1(n46), .A2(IN4[20]), .B1(n13), .B2(IN1[19]), .ZN(n22) );
  AOI22_X1 U18 ( .A1(n48), .A2(IN4[19]), .B1(n12), .B2(IN1[18]), .ZN(n21) );
  NAND2_X1 U19 ( .A1(n22), .A2(n21), .ZN(Y[19]) );
  AOI22_X1 U20 ( .A1(n46), .A2(IN4[21]), .B1(n13), .B2(IN1[20]), .ZN(n24) );
  AOI22_X1 U21 ( .A1(n48), .A2(IN4[20]), .B1(n12), .B2(IN1[19]), .ZN(n23) );
  NAND2_X1 U22 ( .A1(n24), .A2(n23), .ZN(Y[20]) );
  AOI22_X1 U23 ( .A1(n46), .A2(IN4[22]), .B1(n13), .B2(IN1[21]), .ZN(n26) );
  AOI22_X1 U24 ( .A1(n48), .A2(IN4[21]), .B1(n12), .B2(IN1[20]), .ZN(n25) );
  NAND2_X1 U25 ( .A1(n26), .A2(n25), .ZN(Y[21]) );
  AOI22_X1 U26 ( .A1(n46), .A2(IN4[23]), .B1(n13), .B2(IN1[22]), .ZN(n28) );
  AOI22_X1 U27 ( .A1(n48), .A2(IN4[22]), .B1(n12), .B2(IN1[21]), .ZN(n27) );
  NAND2_X1 U28 ( .A1(n28), .A2(n27), .ZN(Y[22]) );
  AOI22_X1 U29 ( .A1(n46), .A2(IN4[24]), .B1(n13), .B2(IN1[23]), .ZN(n30) );
  AOI22_X1 U30 ( .A1(n48), .A2(IN4[23]), .B1(n12), .B2(IN1[22]), .ZN(n29) );
  NAND2_X1 U31 ( .A1(n30), .A2(n29), .ZN(Y[23]) );
  AOI22_X1 U32 ( .A1(n46), .A2(IN4[25]), .B1(n13), .B2(IN1[24]), .ZN(n32) );
  AOI22_X1 U33 ( .A1(n48), .A2(IN4[24]), .B1(n12), .B2(IN1[23]), .ZN(n31) );
  NAND2_X1 U34 ( .A1(n32), .A2(n31), .ZN(Y[24]) );
  AOI22_X1 U35 ( .A1(n46), .A2(IN4[26]), .B1(n13), .B2(IN1[25]), .ZN(n34) );
  AOI22_X1 U36 ( .A1(n48), .A2(IN4[25]), .B1(n12), .B2(IN1[24]), .ZN(n33) );
  NAND2_X1 U37 ( .A1(n34), .A2(n33), .ZN(Y[25]) );
  AOI22_X1 U38 ( .A1(n46), .A2(IN4[27]), .B1(n13), .B2(IN1[26]), .ZN(n36) );
  AOI22_X1 U39 ( .A1(n48), .A2(IN4[26]), .B1(n12), .B2(IN1[25]), .ZN(n35) );
  NAND2_X1 U40 ( .A1(n36), .A2(n35), .ZN(Y[26]) );
  AOI22_X1 U41 ( .A1(n46), .A2(IN4[28]), .B1(n13), .B2(IN1[27]), .ZN(n38) );
  AOI22_X1 U42 ( .A1(n48), .A2(IN4[27]), .B1(n12), .B2(IN1[26]), .ZN(n37) );
  NAND2_X1 U43 ( .A1(n38), .A2(n37), .ZN(Y[27]) );
  AOI22_X1 U44 ( .A1(n46), .A2(IN4[29]), .B1(n13), .B2(IN1[28]), .ZN(n40) );
  AOI22_X1 U45 ( .A1(n48), .A2(IN4[28]), .B1(n12), .B2(IN1[27]), .ZN(n39) );
  NAND2_X1 U46 ( .A1(n40), .A2(n39), .ZN(Y[28]) );
  AOI22_X1 U47 ( .A1(n46), .A2(IN4[30]), .B1(n13), .B2(IN1[29]), .ZN(n42) );
  AOI22_X1 U48 ( .A1(n48), .A2(IN4[29]), .B1(n12), .B2(IN1[28]), .ZN(n41) );
  NAND2_X1 U49 ( .A1(n42), .A2(n41), .ZN(Y[29]) );
  AOI22_X1 U50 ( .A1(n46), .A2(IN4[31]), .B1(n13), .B2(IN1[30]), .ZN(n44) );
  AOI22_X1 U51 ( .A1(n48), .A2(IN4[30]), .B1(n12), .B2(IN1[29]), .ZN(n43) );
  NAND2_X1 U52 ( .A1(n44), .A2(n43), .ZN(Y[30]) );
  AOI22_X1 U53 ( .A1(n46), .A2(IN2[31]), .B1(n13), .B2(IN1[31]), .ZN(n50) );
  AOI22_X1 U54 ( .A1(n48), .A2(IN4[31]), .B1(n12), .B2(IN1[30]), .ZN(n49) );
  NAND2_X1 U55 ( .A1(n50), .A2(n49), .ZN(Y[31]) );
endmodule


module MUX_8to1_N64_7 ( IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, SEL, Y );
  input [63:0] IN0;
  input [63:0] IN1;
  input [63:0] IN2;
  input [63:0] IN3;
  input [63:0] IN4;
  input [63:0] IN5;
  input [63:0] IN6;
  input [63:0] IN7;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n1, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46;

  OAI21_X1 U1 ( .B1(n44), .B2(n43), .A(IN1[18]), .ZN(n1) );
  NAND2_X1 U2 ( .A1(n1), .A2(n18), .ZN(Y[19]) );
  INV_X1 U3 ( .A(n16), .ZN(Y[18]) );
  AND2_X1 U4 ( .A1(n14), .A2(SEL[1]), .ZN(n43) );
  BUF_X1 U5 ( .A(n41), .Z(n12) );
  AND2_X1 U6 ( .A1(SEL[1]), .A2(n13), .ZN(n42) );
  NOR2_X1 U7 ( .A1(n17), .A2(SEL[2]), .ZN(n14) );
  NAND2_X1 U8 ( .A1(n17), .A2(SEL[2]), .ZN(n15) );
  NOR2_X1 U9 ( .A1(SEL[2]), .A2(SEL[0]), .ZN(n13) );
  NOR2_X2 U10 ( .A1(n15), .A2(SEL[1]), .ZN(n44) );
  NOR3_X2 U11 ( .A1(SEL[2]), .A2(SEL[1]), .A3(n17), .ZN(n41) );
  INV_X1 U12 ( .A(SEL[0]), .ZN(n17) );
  OAI21_X1 U13 ( .B1(n42), .B2(n41), .A(IN1[18]), .ZN(n16) );
  AOI22_X1 U14 ( .A1(n42), .A2(IN4[20]), .B1(n41), .B2(IN1[19]), .ZN(n18) );
  AOI22_X1 U15 ( .A1(n42), .A2(IN4[21]), .B1(n41), .B2(IN1[20]), .ZN(n20) );
  AOI22_X1 U16 ( .A1(n44), .A2(IN4[20]), .B1(n43), .B2(IN1[19]), .ZN(n19) );
  NAND2_X1 U17 ( .A1(n20), .A2(n19), .ZN(Y[20]) );
  AOI22_X1 U18 ( .A1(n42), .A2(IN4[22]), .B1(n41), .B2(IN1[21]), .ZN(n22) );
  AOI22_X1 U19 ( .A1(n44), .A2(IN4[21]), .B1(n43), .B2(IN1[20]), .ZN(n21) );
  NAND2_X1 U20 ( .A1(n22), .A2(n21), .ZN(Y[21]) );
  AOI22_X1 U21 ( .A1(n42), .A2(IN4[23]), .B1(n41), .B2(IN1[22]), .ZN(n24) );
  AOI22_X1 U22 ( .A1(n44), .A2(IN4[22]), .B1(n43), .B2(IN1[21]), .ZN(n23) );
  NAND2_X1 U23 ( .A1(n24), .A2(n23), .ZN(Y[22]) );
  AOI22_X1 U24 ( .A1(n42), .A2(IN4[24]), .B1(n41), .B2(IN1[23]), .ZN(n26) );
  AOI22_X1 U25 ( .A1(n44), .A2(IN4[23]), .B1(n43), .B2(IN1[22]), .ZN(n25) );
  NAND2_X1 U26 ( .A1(n26), .A2(n25), .ZN(Y[23]) );
  AOI22_X1 U27 ( .A1(n42), .A2(IN4[25]), .B1(n41), .B2(IN1[24]), .ZN(n28) );
  AOI22_X1 U28 ( .A1(n44), .A2(IN4[24]), .B1(n43), .B2(IN1[23]), .ZN(n27) );
  NAND2_X1 U29 ( .A1(n28), .A2(n27), .ZN(Y[24]) );
  AOI22_X1 U30 ( .A1(n42), .A2(IN4[26]), .B1(n41), .B2(IN1[25]), .ZN(n30) );
  AOI22_X1 U31 ( .A1(n44), .A2(IN4[25]), .B1(n43), .B2(IN1[24]), .ZN(n29) );
  NAND2_X1 U32 ( .A1(n30), .A2(n29), .ZN(Y[25]) );
  AOI22_X1 U33 ( .A1(n42), .A2(IN4[27]), .B1(n41), .B2(IN1[26]), .ZN(n32) );
  AOI22_X1 U34 ( .A1(n44), .A2(IN4[26]), .B1(n43), .B2(IN1[25]), .ZN(n31) );
  NAND2_X1 U35 ( .A1(n32), .A2(n31), .ZN(Y[26]) );
  AOI22_X1 U36 ( .A1(n42), .A2(IN4[28]), .B1(n12), .B2(IN1[27]), .ZN(n34) );
  AOI22_X1 U37 ( .A1(n44), .A2(IN4[27]), .B1(n43), .B2(IN1[26]), .ZN(n33) );
  NAND2_X1 U38 ( .A1(n34), .A2(n33), .ZN(Y[27]) );
  AOI22_X1 U39 ( .A1(n42), .A2(IN4[29]), .B1(n12), .B2(IN1[28]), .ZN(n36) );
  AOI22_X1 U40 ( .A1(n44), .A2(IN4[28]), .B1(n43), .B2(IN1[27]), .ZN(n35) );
  NAND2_X1 U41 ( .A1(n36), .A2(n35), .ZN(Y[28]) );
  AOI22_X1 U42 ( .A1(n42), .A2(IN4[30]), .B1(n12), .B2(IN1[29]), .ZN(n38) );
  AOI22_X1 U43 ( .A1(n44), .A2(IN4[29]), .B1(n43), .B2(IN1[28]), .ZN(n37) );
  NAND2_X1 U44 ( .A1(n38), .A2(n37), .ZN(Y[29]) );
  AOI22_X1 U45 ( .A1(n42), .A2(IN4[31]), .B1(n12), .B2(IN1[30]), .ZN(n40) );
  AOI22_X1 U46 ( .A1(n44), .A2(IN4[30]), .B1(n43), .B2(IN1[29]), .ZN(n39) );
  NAND2_X1 U47 ( .A1(n40), .A2(n39), .ZN(Y[30]) );
  AOI22_X1 U48 ( .A1(n42), .A2(IN2[31]), .B1(n12), .B2(IN1[31]), .ZN(n46) );
  AOI22_X1 U49 ( .A1(n44), .A2(IN4[31]), .B1(n43), .B2(IN1[30]), .ZN(n45) );
  NAND2_X1 U50 ( .A1(n46), .A2(n45), .ZN(Y[31]) );
endmodule


module MUX_8to1_N64_6 ( IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, SEL, Y );
  input [63:0] IN0;
  input [63:0] IN1;
  input [63:0] IN2;
  input [63:0] IN3;
  input [63:0] IN4;
  input [63:0] IN5;
  input [63:0] IN6;
  input [63:0] IN7;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36;

  INV_X1 U1 ( .A(n8), .ZN(Y[20]) );
  AND3_X1 U2 ( .A1(n10), .A2(n9), .A3(SEL[2]), .ZN(n34) );
  NOR3_X2 U3 ( .A1(SEL[2]), .A2(n10), .A3(n9), .ZN(n33) );
  NOR3_X2 U4 ( .A1(SEL[2]), .A2(SEL[1]), .A3(n9), .ZN(n31) );
  NOR3_X2 U5 ( .A1(SEL[2]), .A2(SEL[0]), .A3(n10), .ZN(n32) );
  INV_X1 U6 ( .A(SEL[1]), .ZN(n10) );
  INV_X1 U7 ( .A(SEL[0]), .ZN(n9) );
  OAI21_X1 U8 ( .B1(n32), .B2(n31), .A(IN1[20]), .ZN(n8) );
  OAI21_X1 U9 ( .B1(n34), .B2(n33), .A(IN1[20]), .ZN(n12) );
  AOI22_X1 U10 ( .A1(n32), .A2(IN4[22]), .B1(n31), .B2(IN1[21]), .ZN(n11) );
  NAND2_X1 U11 ( .A1(n12), .A2(n11), .ZN(Y[21]) );
  AOI22_X1 U12 ( .A1(n32), .A2(IN4[23]), .B1(n31), .B2(IN1[22]), .ZN(n14) );
  AOI22_X1 U13 ( .A1(n34), .A2(IN4[22]), .B1(n33), .B2(IN1[21]), .ZN(n13) );
  NAND2_X1 U14 ( .A1(n14), .A2(n13), .ZN(Y[22]) );
  AOI22_X1 U15 ( .A1(n32), .A2(IN4[24]), .B1(n31), .B2(IN1[23]), .ZN(n16) );
  AOI22_X1 U16 ( .A1(n34), .A2(IN4[23]), .B1(n33), .B2(IN1[22]), .ZN(n15) );
  NAND2_X1 U17 ( .A1(n16), .A2(n15), .ZN(Y[23]) );
  AOI22_X1 U18 ( .A1(n32), .A2(IN4[25]), .B1(n31), .B2(IN1[24]), .ZN(n18) );
  AOI22_X1 U19 ( .A1(n34), .A2(IN4[24]), .B1(n33), .B2(IN1[23]), .ZN(n17) );
  NAND2_X1 U20 ( .A1(n18), .A2(n17), .ZN(Y[24]) );
  AOI22_X1 U21 ( .A1(n32), .A2(IN4[26]), .B1(n31), .B2(IN1[25]), .ZN(n20) );
  AOI22_X1 U22 ( .A1(n34), .A2(IN4[25]), .B1(n33), .B2(IN1[24]), .ZN(n19) );
  NAND2_X1 U23 ( .A1(n20), .A2(n19), .ZN(Y[25]) );
  AOI22_X1 U24 ( .A1(n32), .A2(IN4[27]), .B1(n31), .B2(IN1[26]), .ZN(n22) );
  AOI22_X1 U25 ( .A1(n34), .A2(IN4[26]), .B1(n33), .B2(IN1[25]), .ZN(n21) );
  NAND2_X1 U26 ( .A1(n22), .A2(n21), .ZN(Y[26]) );
  AOI22_X1 U27 ( .A1(n32), .A2(IN4[28]), .B1(n31), .B2(IN1[27]), .ZN(n24) );
  AOI22_X1 U28 ( .A1(n34), .A2(IN4[27]), .B1(n33), .B2(IN1[26]), .ZN(n23) );
  NAND2_X1 U29 ( .A1(n24), .A2(n23), .ZN(Y[27]) );
  AOI22_X1 U30 ( .A1(n32), .A2(IN4[29]), .B1(n31), .B2(IN1[28]), .ZN(n26) );
  AOI22_X1 U31 ( .A1(n34), .A2(IN4[28]), .B1(n33), .B2(IN1[27]), .ZN(n25) );
  NAND2_X1 U32 ( .A1(n26), .A2(n25), .ZN(Y[28]) );
  AOI22_X1 U33 ( .A1(n32), .A2(IN4[30]), .B1(n31), .B2(IN1[29]), .ZN(n28) );
  AOI22_X1 U34 ( .A1(n34), .A2(IN4[29]), .B1(n33), .B2(IN1[28]), .ZN(n27) );
  NAND2_X1 U35 ( .A1(n28), .A2(n27), .ZN(Y[29]) );
  AOI22_X1 U36 ( .A1(n32), .A2(IN4[31]), .B1(n31), .B2(IN1[30]), .ZN(n30) );
  AOI22_X1 U37 ( .A1(n34), .A2(IN4[30]), .B1(n33), .B2(IN1[29]), .ZN(n29) );
  NAND2_X1 U38 ( .A1(n30), .A2(n29), .ZN(Y[30]) );
  AOI22_X1 U39 ( .A1(n32), .A2(IN2[31]), .B1(n31), .B2(IN1[31]), .ZN(n36) );
  AOI22_X1 U40 ( .A1(n34), .A2(IN4[31]), .B1(n33), .B2(IN1[30]), .ZN(n35) );
  NAND2_X1 U41 ( .A1(n36), .A2(n35), .ZN(Y[31]) );
endmodule


module MUX_8to1_N64_5 ( IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, SEL, Y );
  input [63:0] IN0;
  input [63:0] IN1;
  input [63:0] IN2;
  input [63:0] IN3;
  input [63:0] IN4;
  input [63:0] IN5;
  input [63:0] IN6;
  input [63:0] IN7;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32;

  INV_X1 U1 ( .A(n8), .ZN(Y[22]) );
  AND3_X1 U2 ( .A1(n10), .A2(n9), .A3(SEL[2]), .ZN(n30) );
  NOR3_X2 U3 ( .A1(SEL[2]), .A2(n10), .A3(n9), .ZN(n29) );
  NOR3_X2 U4 ( .A1(SEL[2]), .A2(SEL[1]), .A3(n9), .ZN(n27) );
  NOR3_X2 U5 ( .A1(SEL[2]), .A2(SEL[0]), .A3(n10), .ZN(n28) );
  INV_X1 U6 ( .A(SEL[1]), .ZN(n10) );
  INV_X1 U7 ( .A(SEL[0]), .ZN(n9) );
  OAI21_X1 U8 ( .B1(n28), .B2(n27), .A(IN1[22]), .ZN(n8) );
  OAI21_X1 U9 ( .B1(n30), .B2(n29), .A(IN1[22]), .ZN(n12) );
  AOI22_X1 U10 ( .A1(n28), .A2(IN4[24]), .B1(n27), .B2(IN1[23]), .ZN(n11) );
  NAND2_X1 U11 ( .A1(n12), .A2(n11), .ZN(Y[23]) );
  AOI22_X1 U12 ( .A1(n28), .A2(IN4[25]), .B1(n27), .B2(IN1[24]), .ZN(n14) );
  AOI22_X1 U13 ( .A1(n30), .A2(IN4[24]), .B1(n29), .B2(IN1[23]), .ZN(n13) );
  NAND2_X1 U14 ( .A1(n14), .A2(n13), .ZN(Y[24]) );
  AOI22_X1 U15 ( .A1(n28), .A2(IN4[26]), .B1(n27), .B2(IN1[25]), .ZN(n16) );
  AOI22_X1 U16 ( .A1(n30), .A2(IN4[25]), .B1(n29), .B2(IN1[24]), .ZN(n15) );
  NAND2_X1 U17 ( .A1(n16), .A2(n15), .ZN(Y[25]) );
  AOI22_X1 U18 ( .A1(n28), .A2(IN4[27]), .B1(n27), .B2(IN1[26]), .ZN(n18) );
  AOI22_X1 U19 ( .A1(n30), .A2(IN4[26]), .B1(n29), .B2(IN1[25]), .ZN(n17) );
  NAND2_X1 U20 ( .A1(n18), .A2(n17), .ZN(Y[26]) );
  AOI22_X1 U21 ( .A1(n28), .A2(IN4[28]), .B1(n27), .B2(IN1[27]), .ZN(n20) );
  AOI22_X1 U22 ( .A1(n30), .A2(IN4[27]), .B1(n29), .B2(IN1[26]), .ZN(n19) );
  NAND2_X1 U23 ( .A1(n20), .A2(n19), .ZN(Y[27]) );
  AOI22_X1 U24 ( .A1(n28), .A2(IN4[29]), .B1(n27), .B2(IN1[28]), .ZN(n22) );
  AOI22_X1 U25 ( .A1(n30), .A2(IN4[28]), .B1(n29), .B2(IN1[27]), .ZN(n21) );
  NAND2_X1 U26 ( .A1(n22), .A2(n21), .ZN(Y[28]) );
  AOI22_X1 U27 ( .A1(n28), .A2(IN4[30]), .B1(n27), .B2(IN1[29]), .ZN(n24) );
  AOI22_X1 U28 ( .A1(n30), .A2(IN4[29]), .B1(n29), .B2(IN1[28]), .ZN(n23) );
  NAND2_X1 U29 ( .A1(n24), .A2(n23), .ZN(Y[29]) );
  AOI22_X1 U30 ( .A1(n28), .A2(IN4[31]), .B1(n27), .B2(IN1[30]), .ZN(n26) );
  AOI22_X1 U31 ( .A1(n30), .A2(IN4[30]), .B1(n29), .B2(IN1[29]), .ZN(n25) );
  NAND2_X1 U32 ( .A1(n26), .A2(n25), .ZN(Y[30]) );
  AOI22_X1 U33 ( .A1(n28), .A2(IN2[31]), .B1(n27), .B2(IN1[31]), .ZN(n32) );
  AOI22_X1 U34 ( .A1(n30), .A2(IN4[31]), .B1(n29), .B2(IN1[30]), .ZN(n31) );
  NAND2_X1 U35 ( .A1(n32), .A2(n31), .ZN(Y[31]) );
endmodule


module MUX_8to1_N64_4 ( IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, SEL, Y );
  input [63:0] IN0;
  input [63:0] IN1;
  input [63:0] IN2;
  input [63:0] IN3;
  input [63:0] IN4;
  input [63:0] IN5;
  input [63:0] IN6;
  input [63:0] IN7;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27;

  AND3_X1 U1 ( .A1(n9), .A2(n8), .A3(SEL[2]), .ZN(n25) );
  NOR3_X2 U2 ( .A1(SEL[2]), .A2(SEL[1]), .A3(n8), .ZN(n22) );
  NOR3_X2 U3 ( .A1(SEL[2]), .A2(SEL[0]), .A3(n9), .ZN(n23) );
  INV_X1 U4 ( .A(SEL[1]), .ZN(n9) );
  INV_X1 U5 ( .A(SEL[0]), .ZN(n8) );
  OAI21_X1 U6 ( .B1(n23), .B2(n22), .A(IN1[24]), .ZN(n7) );
  INV_X1 U7 ( .A(n7), .ZN(Y[24]) );
  NOR3_X1 U8 ( .A1(SEL[2]), .A2(n9), .A3(n8), .ZN(n24) );
  OAI21_X1 U9 ( .B1(n25), .B2(n24), .A(IN1[24]), .ZN(n11) );
  AOI22_X1 U10 ( .A1(n23), .A2(IN4[26]), .B1(n22), .B2(IN1[25]), .ZN(n10) );
  NAND2_X1 U11 ( .A1(n11), .A2(n10), .ZN(Y[25]) );
  AOI22_X1 U12 ( .A1(n23), .A2(IN4[27]), .B1(n22), .B2(IN1[26]), .ZN(n13) );
  AOI22_X1 U13 ( .A1(n25), .A2(IN4[26]), .B1(n24), .B2(IN1[25]), .ZN(n12) );
  NAND2_X1 U14 ( .A1(n13), .A2(n12), .ZN(Y[26]) );
  AOI22_X1 U15 ( .A1(n23), .A2(IN4[28]), .B1(n22), .B2(IN1[27]), .ZN(n15) );
  AOI22_X1 U16 ( .A1(n25), .A2(IN4[27]), .B1(n24), .B2(IN1[26]), .ZN(n14) );
  NAND2_X1 U17 ( .A1(n15), .A2(n14), .ZN(Y[27]) );
  AOI22_X1 U18 ( .A1(n23), .A2(IN4[29]), .B1(n22), .B2(IN1[28]), .ZN(n17) );
  AOI22_X1 U19 ( .A1(n25), .A2(IN4[28]), .B1(n24), .B2(IN1[27]), .ZN(n16) );
  NAND2_X1 U20 ( .A1(n17), .A2(n16), .ZN(Y[28]) );
  AOI22_X1 U21 ( .A1(n23), .A2(IN4[30]), .B1(n22), .B2(IN1[29]), .ZN(n19) );
  AOI22_X1 U22 ( .A1(n25), .A2(IN4[29]), .B1(n24), .B2(IN1[28]), .ZN(n18) );
  NAND2_X1 U23 ( .A1(n19), .A2(n18), .ZN(Y[29]) );
  AOI22_X1 U24 ( .A1(n23), .A2(IN4[31]), .B1(n22), .B2(IN1[30]), .ZN(n21) );
  AOI22_X1 U25 ( .A1(n25), .A2(IN4[30]), .B1(n24), .B2(IN1[29]), .ZN(n20) );
  NAND2_X1 U26 ( .A1(n21), .A2(n20), .ZN(Y[30]) );
  AOI22_X1 U27 ( .A1(n23), .A2(IN2[31]), .B1(n22), .B2(IN1[31]), .ZN(n27) );
  AOI22_X1 U28 ( .A1(n25), .A2(IN4[31]), .B1(n24), .B2(IN1[30]), .ZN(n26) );
  NAND2_X1 U29 ( .A1(n27), .A2(n26), .ZN(Y[31]) );
endmodule


module MUX_8to1_N64_3 ( IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, SEL, Y );
  input [63:0] IN0;
  input [63:0] IN1;
  input [63:0] IN2;
  input [63:0] IN3;
  input [63:0] IN4;
  input [63:0] IN5;
  input [63:0] IN6;
  input [63:0] IN7;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n1, n2, n3, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28;

  BUF_X1 U1 ( .A(SEL[1]), .Z(n1) );
  BUF_X2 U2 ( .A(n23), .Z(n2) );
  BUF_X1 U3 ( .A(n26), .Z(n3) );
  NOR2_X1 U4 ( .A1(n11), .A2(n1), .ZN(n26) );
  AND2_X2 U5 ( .A1(n12), .A2(n1), .ZN(n25) );
  BUF_X1 U6 ( .A(SEL[0]), .Z(n9) );
  NOR3_X1 U7 ( .A1(SEL[2]), .A2(SEL[1]), .A3(n14), .ZN(n23) );
  AND2_X2 U8 ( .A1(n10), .A2(n1), .ZN(n24) );
  NOR2_X1 U9 ( .A1(n14), .A2(SEL[2]), .ZN(n12) );
  NAND2_X1 U10 ( .A1(n14), .A2(SEL[2]), .ZN(n11) );
  NOR2_X1 U11 ( .A1(SEL[2]), .A2(n9), .ZN(n10) );
  INV_X1 U12 ( .A(SEL[0]), .ZN(n14) );
  OAI21_X1 U13 ( .B1(n24), .B2(n2), .A(IN1[26]), .ZN(n13) );
  INV_X1 U14 ( .A(n13), .ZN(Y[26]) );
  OAI21_X1 U15 ( .B1(n26), .B2(n25), .A(IN1[26]), .ZN(n16) );
  AOI22_X1 U16 ( .A1(n24), .A2(IN4[28]), .B1(n2), .B2(IN1[27]), .ZN(n15) );
  NAND2_X1 U17 ( .A1(n16), .A2(n15), .ZN(Y[27]) );
  AOI22_X1 U18 ( .A1(n24), .A2(IN4[29]), .B1(n2), .B2(IN1[28]), .ZN(n18) );
  AOI22_X1 U19 ( .A1(n26), .A2(IN4[28]), .B1(n25), .B2(IN1[27]), .ZN(n17) );
  NAND2_X1 U20 ( .A1(n18), .A2(n17), .ZN(Y[28]) );
  AOI22_X1 U21 ( .A1(n24), .A2(IN4[30]), .B1(n2), .B2(IN1[29]), .ZN(n20) );
  AOI22_X1 U22 ( .A1(n26), .A2(IN4[29]), .B1(n25), .B2(IN1[28]), .ZN(n19) );
  NAND2_X1 U23 ( .A1(n20), .A2(n19), .ZN(Y[29]) );
  AOI22_X1 U24 ( .A1(n24), .A2(IN4[31]), .B1(n2), .B2(IN1[30]), .ZN(n22) );
  AOI22_X1 U25 ( .A1(n3), .A2(IN4[30]), .B1(n25), .B2(IN1[29]), .ZN(n21) );
  NAND2_X1 U26 ( .A1(n22), .A2(n21), .ZN(Y[30]) );
  AOI22_X1 U27 ( .A1(n24), .A2(IN2[31]), .B1(n2), .B2(IN1[31]), .ZN(n28) );
  AOI22_X1 U28 ( .A1(n3), .A2(IN4[31]), .B1(n25), .B2(IN1[30]), .ZN(n27) );
  NAND2_X1 U29 ( .A1(n28), .A2(n27), .ZN(Y[31]) );
endmodule


module MUX_8to1_N64_2 ( IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, SEL, Y );
  input [63:0] IN0;
  input [63:0] IN1;
  input [63:0] IN2;
  input [63:0] IN3;
  input [63:0] IN4;
  input [63:0] IN5;
  input [63:0] IN6;
  input [63:0] IN7;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17;

  INV_X1 U1 ( .A(SEL[1]), .ZN(n7) );
  NOR3_X1 U2 ( .A1(SEL[2]), .A2(SEL[0]), .A3(n7), .ZN(n13) );
  INV_X1 U3 ( .A(SEL[0]), .ZN(n6) );
  NOR3_X1 U4 ( .A1(SEL[2]), .A2(SEL[1]), .A3(n6), .ZN(n12) );
  OAI21_X1 U5 ( .B1(n13), .B2(n12), .A(IN1[28]), .ZN(n5) );
  INV_X1 U6 ( .A(n5), .ZN(Y[28]) );
  AND3_X1 U7 ( .A1(n7), .A2(n6), .A3(SEL[2]), .ZN(n15) );
  NOR3_X1 U8 ( .A1(SEL[2]), .A2(n7), .A3(n6), .ZN(n14) );
  OAI21_X1 U9 ( .B1(n15), .B2(n14), .A(IN1[28]), .ZN(n9) );
  AOI22_X1 U10 ( .A1(n13), .A2(IN4[30]), .B1(n12), .B2(IN1[29]), .ZN(n8) );
  NAND2_X1 U11 ( .A1(n9), .A2(n8), .ZN(Y[29]) );
  AOI22_X1 U12 ( .A1(n13), .A2(IN4[31]), .B1(n12), .B2(IN1[30]), .ZN(n11) );
  AOI22_X1 U13 ( .A1(n15), .A2(IN4[30]), .B1(n14), .B2(IN1[29]), .ZN(n10) );
  NAND2_X1 U14 ( .A1(n11), .A2(n10), .ZN(Y[30]) );
  AOI22_X1 U15 ( .A1(n13), .A2(IN2[31]), .B1(n12), .B2(IN1[31]), .ZN(n17) );
  AOI22_X1 U16 ( .A1(n15), .A2(IN4[31]), .B1(n14), .B2(IN1[30]), .ZN(n16) );
  NAND2_X1 U17 ( .A1(n17), .A2(n16), .ZN(Y[31]) );
endmodule


module MUX_8to1_N64_1 ( IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, SEL, Y );
  input [63:0] IN0;
  input [63:0] IN1;
  input [63:0] IN2;
  input [63:0] IN3;
  input [63:0] IN4;
  input [63:0] IN5;
  input [63:0] IN6;
  input [63:0] IN7;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n3, n4, n5, n6, n7, n8, n9;

  INV_X1 U1 ( .A(SEL[2]), .ZN(n4) );
  OAI211_X1 U2 ( .C1(SEL[1]), .C2(SEL[0]), .A(IN1[30]), .B(n4), .ZN(n3) );
  AOI21_X1 U3 ( .B1(SEL[1]), .B2(SEL[0]), .A(n3), .ZN(Y[30]) );
  NOR2_X1 U4 ( .A1(SEL[0]), .A2(n4), .ZN(n6) );
  INV_X1 U5 ( .A(SEL[0]), .ZN(n7) );
  NOR2_X1 U6 ( .A1(SEL[2]), .A2(n7), .ZN(n5) );
  AOI22_X1 U7 ( .A1(IN1[30]), .A2(n6), .B1(IN1[31]), .B2(n5), .ZN(n9) );
  OAI221_X1 U8 ( .B1(SEL[0]), .B2(IN2[31]), .C1(n7), .C2(IN1[30]), .A(SEL[1]), 
        .ZN(n8) );
  OAI22_X1 U9 ( .A1(SEL[1]), .A2(n9), .B1(SEL[2]), .B2(n8), .ZN(Y[31]) );
endmodule


module booth_encoder_0 ( \input , \output  );
  input [1:-1] \input ;
  output [2:0] \output ;
  wire   n1, n2;

  NOR2_X1 U1 ( .A1(n2), .A2(\input [0]), .ZN(\output [2]) );
  INV_X1 U2 ( .A(\input [1]), .ZN(n2) );
  NOR2_X1 U3 ( .A1(n1), .A2(\input [1]), .ZN(\output [0]) );
  INV_X1 U4 ( .A(\input [0]), .ZN(n1) );
  NOR2_X1 U5 ( .A1(n2), .A2(n1), .ZN(\output [1]) );
endmodule


module booth_encoder_15 ( \input , \output  );
  input [1:-1] \input ;
  output [2:0] \output ;
  wire   n1, n2, n3;

  NOR2_X1 U1 ( .A1(\input [-1]), .A2(\input [0]), .ZN(n3) );
  AND2_X1 U2 ( .A1(\input [1]), .A2(n3), .ZN(\output [2]) );
  NOR2_X1 U3 ( .A1(n3), .A2(\input [1]), .ZN(\output [0]) );
  NAND2_X1 U4 ( .A1(\input [-1]), .A2(\input [0]), .ZN(n1) );
  NAND2_X1 U5 ( .A1(n1), .A2(\input [1]), .ZN(n2) );
  OAI22_X1 U6 ( .A1(n2), .A2(n3), .B1(n1), .B2(\input [1]), .ZN(\output [1])
         );
endmodule


module booth_encoder_14 ( \input , \output  );
  input [1:-1] \input ;
  output [2:0] \output ;
  wire   n1, n2, n3;

  NOR2_X1 U1 ( .A1(\input [0]), .A2(\input [-1]), .ZN(n3) );
  AND2_X1 U2 ( .A1(n3), .A2(\input [1]), .ZN(\output [2]) );
  NOR2_X1 U3 ( .A1(n3), .A2(\input [1]), .ZN(\output [0]) );
  NAND2_X1 U4 ( .A1(\input [-1]), .A2(\input [0]), .ZN(n1) );
  NAND2_X1 U5 ( .A1(\input [1]), .A2(n1), .ZN(n2) );
  OAI22_X1 U6 ( .A1(n3), .A2(n2), .B1(\input [1]), .B2(n1), .ZN(\output [1])
         );
endmodule


module booth_encoder_13 ( \input , \output  );
  input [1:-1] \input ;
  output [2:0] \output ;
  wire   n1, n2, n3;

  NOR2_X1 U1 ( .A1(\input [0]), .A2(\input [-1]), .ZN(n3) );
  AND2_X1 U2 ( .A1(n3), .A2(\input [1]), .ZN(\output [2]) );
  NOR2_X1 U3 ( .A1(n3), .A2(\input [1]), .ZN(\output [0]) );
  NAND2_X1 U4 ( .A1(\input [0]), .A2(\input [-1]), .ZN(n1) );
  NAND2_X1 U5 ( .A1(\input [1]), .A2(n1), .ZN(n2) );
  OAI22_X1 U6 ( .A1(n3), .A2(n2), .B1(\input [1]), .B2(n1), .ZN(\output [1])
         );
endmodule


module booth_encoder_12 ( \input , \output  );
  input [1:-1] \input ;
  output [2:0] \output ;
  wire   n2, n3, n4;

  AND2_X1 U1 ( .A1(n4), .A2(\input [1]), .ZN(\output [2]) );
  NOR2_X1 U2 ( .A1(\input [0]), .A2(\input [-1]), .ZN(n4) );
  NOR2_X1 U3 ( .A1(n4), .A2(\input [1]), .ZN(\output [0]) );
  NAND2_X1 U4 ( .A1(\input [0]), .A2(\input [-1]), .ZN(n2) );
  NAND2_X1 U5 ( .A1(\input [1]), .A2(n2), .ZN(n3) );
  OAI22_X1 U6 ( .A1(n4), .A2(n3), .B1(\input [1]), .B2(n2), .ZN(\output [1])
         );
endmodule


module booth_encoder_11 ( \input , \output  );
  input [1:-1] \input ;
  output [2:0] \output ;
  wire   n2, n3, n4;

  OAI22_X1 U1 ( .A1(n2), .A2(n4), .B1(n3), .B2(\input [1]), .ZN(\output [1])
         );
  NAND2_X1 U2 ( .A1(n3), .A2(\input [1]), .ZN(n2) );
  AND2_X1 U3 ( .A1(\input [1]), .A2(n4), .ZN(\output [2]) );
  NOR2_X1 U4 ( .A1(\input [0]), .A2(\input [-1]), .ZN(n4) );
  NOR2_X1 U5 ( .A1(n4), .A2(\input [1]), .ZN(\output [0]) );
  NAND2_X1 U6 ( .A1(\input [0]), .A2(\input [-1]), .ZN(n3) );
endmodule


module booth_encoder_10 ( \input , \output  );
  input [1:-1] \input ;
  output [2:0] \output ;
  wire   n1, n2, n3;

  AND2_X1 U1 ( .A1(n3), .A2(\input [1]), .ZN(\output [2]) );
  NOR2_X1 U2 ( .A1(\input [0]), .A2(\input [-1]), .ZN(n3) );
  NOR2_X1 U3 ( .A1(n3), .A2(\input [1]), .ZN(\output [0]) );
  NAND2_X1 U4 ( .A1(\input [0]), .A2(\input [-1]), .ZN(n1) );
  NAND2_X1 U5 ( .A1(\input [1]), .A2(n1), .ZN(n2) );
  OAI22_X1 U6 ( .A1(n3), .A2(n2), .B1(\input [1]), .B2(n1), .ZN(\output [1])
         );
endmodule


module booth_encoder_9 ( \input , \output  );
  input [1:-1] \input ;
  output [2:0] \output ;
  wire   n1, n2, n3;

  AND2_X1 U1 ( .A1(n3), .A2(\input [1]), .ZN(\output [2]) );
  NOR2_X1 U2 ( .A1(\input [0]), .A2(\input [-1]), .ZN(n3) );
  NOR2_X1 U3 ( .A1(n3), .A2(\input [1]), .ZN(\output [0]) );
  NAND2_X1 U4 ( .A1(\input [0]), .A2(\input [-1]), .ZN(n1) );
  NAND2_X1 U5 ( .A1(\input [1]), .A2(n1), .ZN(n2) );
  OAI22_X1 U6 ( .A1(n3), .A2(n2), .B1(\input [1]), .B2(n1), .ZN(\output [1])
         );
endmodule


module booth_encoder_8 ( \input , \output  );
  input [1:-1] \input ;
  output [2:0] \output ;
  wire   n1, n2, n3;

  AND2_X1 U1 ( .A1(n3), .A2(\input [1]), .ZN(\output [2]) );
  NOR2_X1 U2 ( .A1(\input [0]), .A2(\input [-1]), .ZN(n3) );
  NOR2_X1 U3 ( .A1(n3), .A2(\input [1]), .ZN(\output [0]) );
  NAND2_X1 U4 ( .A1(\input [0]), .A2(\input [-1]), .ZN(n1) );
  NAND2_X1 U5 ( .A1(\input [1]), .A2(n1), .ZN(n2) );
  OAI22_X1 U6 ( .A1(n3), .A2(n2), .B1(\input [1]), .B2(n1), .ZN(\output [1])
         );
endmodule


module booth_encoder_7 ( \input , \output  );
  input [1:-1] \input ;
  output [2:0] \output ;
  wire   n1, n2, n3;

  AND2_X1 U1 ( .A1(n3), .A2(\input [1]), .ZN(\output [2]) );
  NOR2_X1 U2 ( .A1(\input [0]), .A2(\input [-1]), .ZN(n3) );
  NOR2_X1 U3 ( .A1(n3), .A2(\input [1]), .ZN(\output [0]) );
  NAND2_X1 U4 ( .A1(\input [0]), .A2(\input [-1]), .ZN(n1) );
  NAND2_X1 U5 ( .A1(\input [1]), .A2(n1), .ZN(n2) );
  OAI22_X1 U6 ( .A1(n3), .A2(n2), .B1(\input [1]), .B2(n1), .ZN(\output [1])
         );
endmodule


module booth_encoder_6 ( \input , \output  );
  input [1:-1] \input ;
  output [2:0] \output ;
  wire   n1, n2, n3;

  AND2_X1 U1 ( .A1(n3), .A2(\input [1]), .ZN(\output [2]) );
  NOR2_X1 U2 ( .A1(\input [0]), .A2(\input [-1]), .ZN(n3) );
  NOR2_X1 U3 ( .A1(n3), .A2(\input [1]), .ZN(\output [0]) );
  NAND2_X1 U4 ( .A1(\input [0]), .A2(\input [-1]), .ZN(n1) );
  NAND2_X1 U5 ( .A1(\input [1]), .A2(n1), .ZN(n2) );
  OAI22_X1 U6 ( .A1(n3), .A2(n2), .B1(\input [1]), .B2(n1), .ZN(\output [1])
         );
endmodule


module booth_encoder_5 ( \input , \output  );
  input [1:-1] \input ;
  output [2:0] \output ;
  wire   n1, n2, n3;

  AND2_X1 U1 ( .A1(n3), .A2(\input [1]), .ZN(\output [2]) );
  NOR2_X1 U2 ( .A1(\input [0]), .A2(\input [-1]), .ZN(n3) );
  NOR2_X1 U3 ( .A1(n3), .A2(\input [1]), .ZN(\output [0]) );
  NAND2_X1 U4 ( .A1(\input [0]), .A2(\input [-1]), .ZN(n1) );
  NAND2_X1 U5 ( .A1(\input [1]), .A2(n1), .ZN(n2) );
  OAI22_X1 U6 ( .A1(n3), .A2(n2), .B1(\input [1]), .B2(n1), .ZN(\output [1])
         );
endmodule


module booth_encoder_4 ( \input , \output  );
  input [1:-1] \input ;
  output [2:0] \output ;
  wire   n2, n3, n4;

  AND2_X1 U1 ( .A1(n4), .A2(\input [1]), .ZN(\output [2]) );
  NOR2_X1 U2 ( .A1(\input [0]), .A2(\input [-1]), .ZN(n4) );
  NOR2_X1 U3 ( .A1(n4), .A2(\input [1]), .ZN(\output [0]) );
  NAND2_X1 U4 ( .A1(\input [0]), .A2(\input [-1]), .ZN(n2) );
  NAND2_X1 U5 ( .A1(\input [1]), .A2(n2), .ZN(n3) );
  OAI22_X1 U6 ( .A1(n4), .A2(n3), .B1(\input [1]), .B2(n2), .ZN(\output [1])
         );
endmodule


module booth_encoder_3 ( \input , \output  );
  input [1:-1] \input ;
  output [2:0] \output ;
  wire   n2, n3, n4;

  AND2_X1 U1 ( .A1(n4), .A2(\input [1]), .ZN(\output [2]) );
  NOR2_X1 U2 ( .A1(\input [0]), .A2(\input [-1]), .ZN(n4) );
  NOR2_X1 U3 ( .A1(n4), .A2(\input [1]), .ZN(\output [0]) );
  NAND2_X1 U4 ( .A1(\input [0]), .A2(\input [-1]), .ZN(n2) );
  NAND2_X1 U5 ( .A1(\input [1]), .A2(n2), .ZN(n3) );
  OAI22_X1 U6 ( .A1(n3), .A2(n4), .B1(\input [1]), .B2(n2), .ZN(\output [1])
         );
endmodule


module booth_encoder_2 ( \input , \output  );
  input [1:-1] \input ;
  output [2:0] \output ;
  wire   n1, n2, n3;

  NOR2_X1 U1 ( .A1(\input [0]), .A2(\input [-1]), .ZN(n3) );
  AND2_X1 U2 ( .A1(n3), .A2(\input [1]), .ZN(\output [2]) );
  NOR2_X1 U3 ( .A1(n3), .A2(\input [1]), .ZN(\output [0]) );
  NAND2_X1 U4 ( .A1(\input [0]), .A2(\input [-1]), .ZN(n1) );
  NAND2_X1 U5 ( .A1(\input [1]), .A2(n1), .ZN(n2) );
  OAI22_X1 U6 ( .A1(n3), .A2(n2), .B1(\input [1]), .B2(n1), .ZN(\output [1])
         );
endmodule


module booth_encoder_1 ( \input , \output  );
  input [1:-1] \input ;
  output [2:0] \output ;
  wire   n1, n2, n3;

  NOR2_X1 U1 ( .A1(\input [0]), .A2(\input [-1]), .ZN(n3) );
  AND2_X1 U2 ( .A1(n3), .A2(\input [1]), .ZN(\output [2]) );
  NOR2_X1 U3 ( .A1(n3), .A2(\input [1]), .ZN(\output [0]) );
  NAND2_X1 U4 ( .A1(\input [0]), .A2(\input [-1]), .ZN(n1) );
  NAND2_X1 U5 ( .A1(\input [1]), .A2(n1), .ZN(n2) );
  OAI22_X1 U6 ( .A1(n3), .A2(n2), .B1(\input [1]), .B2(n1), .ZN(\output [1])
         );
endmodule


module SNPS_CLOCK_GATE_HIGH_boothmul_4stage_N32_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18800, net18802, net18804, net18805, net18808, net18811;
  assign net18800 = EN;
  assign net18802 = CLK;
  assign ENCLK = net18804;
  assign net18811 = TE;

  DLL_X1 latch ( .D(net18805), .GN(net18802), .Q(net18808) );
  AND2_X1 main_gate ( .A1(net18808), .A2(net18802), .ZN(net18804) );
  OR2_X1 test_or ( .A1(net18800), .A2(net18811), .ZN(net18805) );
endmodule


module SNPS_CLOCK_GATE_HIGH_boothmul_4stage_N32_3 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18800, net18802, net18804, net18805, net18808, net18811;
  assign net18800 = EN;
  assign net18802 = CLK;
  assign ENCLK = net18804;
  assign net18811 = TE;

  DLL_X1 latch ( .D(net18805), .GN(net18802), .Q(net18808) );
  AND2_X1 main_gate ( .A1(net18808), .A2(net18802), .ZN(net18804) );
  OR2_X1 test_or ( .A1(net18800), .A2(net18811), .ZN(net18805) );
endmodule


module SNPS_CLOCK_GATE_HIGH_boothmul_4stage_N32_1 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18800, net18802, net18804, net18805, net18808, net18811;
  assign net18800 = EN;
  assign net18802 = CLK;
  assign ENCLK = net18804;
  assign net18811 = TE;

  DLL_X1 latch ( .D(net18805), .GN(net18802), .Q(net18808) );
  AND2_X1 main_gate ( .A1(net18808), .A2(net18802), .ZN(net18804) );
  OR2_X1 test_or ( .A1(net18800), .A2(net18811), .ZN(net18805) );
endmodule


module boothmul_4stage_N32 ( A, B, EN, CLK, RST, P );
  input [31:0] A;
  input [31:0] B;
  output [63:0] P;
  input EN, CLK, RST;
  wire   \add_out_s2[7][31] , \add_out_s2[7][30] , \add_out_s2[7][29] ,
         \add_out_s2[7][27] , \add_out_s2[7][26] , \add_out_s2[7][25] ,
         \add_out_s2[7][24] , \add_out_s2[7][23] , \add_out_s2[7][22] ,
         \add_out_s2[7][21] , \add_out_s2[7][20] , \add_out_s2[7][19] ,
         \add_out_s2[7][18] , \add_out_s2[7][17] , \add_out_s2[7][16] ,
         \add_out_s2[7][15] , \add_out_s2[7][14] , \add_out_s2[7][13] ,
         \add_out_s2[7][12] , \add_out_s2[7][11] , \add_out_s2[7][10] ,
         \add_out_s2[7][9] , \add_out_s2[7][8] , \add_out_s2[7][7] ,
         \add_out_s2[7][6] , \add_out_s2[7][5] , \add_out_s2[7][4] ,
         \add_out_s2[7][3] , \add_out_s2[7][2] , \add_out_s2[7][1] ,
         \add_out_s2[7][0] , \add_out_s2[6][31] , \add_out_s2[6][30] ,
         \add_out_s2[6][29] , \add_out_s2[6][28] , \add_out_s2[6][27] ,
         \add_out_s2[6][26] , \add_out_s2[6][25] , \add_out_s2[6][24] ,
         \add_out_s2[6][23] , \add_out_s2[6][22] , \add_out_s2[6][21] ,
         \add_out_s2[6][20] , \add_out_s2[6][19] , \add_out_s2[6][18] ,
         \add_out_s2[6][17] , \add_out_s2[6][16] , \add_out_s2[6][15] ,
         \add_out_s2[6][14] , \add_out_s2[6][13] , \add_out_s2[6][12] ,
         \add_out_s2[6][11] , \add_out_s2[6][10] , \add_out_s2[6][9] ,
         \add_out_s2[6][8] , \add_out_s2[6][7] , \add_out_s2[6][6] ,
         \add_out_s2[6][5] , \add_out_s2[6][4] , \add_out_s2[6][3] ,
         \add_out_s2[6][2] , \add_out_s2[6][1] , \add_out_s2[6][0] ,
         \add_out_s2[5][31] , \add_out_s2[5][30] , \add_out_s2[5][29] ,
         \add_out_s2[5][28] , \add_out_s2[5][27] , \add_out_s2[5][26] ,
         \add_out_s2[5][25] , \add_out_s2[5][24] , \add_out_s2[5][23] ,
         \add_out_s2[5][22] , \add_out_s2[5][21] , \add_out_s2[5][19] ,
         \add_out_s2[5][18] , \add_out_s2[5][17] , \add_out_s2[5][16] ,
         \add_out_s2[5][15] , \add_out_s2[5][14] , \add_out_s2[5][13] ,
         \add_out_s2[5][12] , \add_out_s2[5][11] , \add_out_s2[5][10] ,
         \add_out_s2[5][9] , \add_out_s2[5][8] , \add_out_s2[5][7] ,
         \add_out_s2[5][6] , \add_out_s2[5][5] , \add_out_s2[5][4] ,
         \add_out_s2[5][3] , \add_out_s2[5][2] , \add_out_s2[5][1] ,
         \add_out_s2[5][0] , \add_out_s2[4][31] , \add_out_s2[4][30] ,
         \add_out_s2[4][29] , \add_out_s2[4][28] , \add_out_s2[4][27] ,
         \add_out_s2[4][26] , \add_out_s2[4][25] , \add_out_s2[4][24] ,
         \add_out_s2[4][23] , \add_out_s2[4][22] , \add_out_s2[4][21] ,
         \add_out_s2[4][20] , \add_out_s2[4][19] , \add_out_s2[4][18] ,
         \add_out_s2[4][17] , \add_out_s2[4][16] , \add_out_s2[4][15] ,
         \add_out_s2[4][14] , \add_out_s2[4][13] , \add_out_s2[4][12] ,
         \add_out_s2[4][11] , \add_out_s2[4][10] , \add_out_s2[4][9] ,
         \add_out_s2[4][8] , \add_out_s2[4][7] , \add_out_s2[4][6] ,
         \add_out_s2[4][5] , \add_out_s2[4][4] , \add_out_s2[4][3] ,
         \add_out_s2[4][2] , \add_out_s2[4][1] , \add_out_s2[4][0] ,
         \add_out_s3[12][31] , \add_out_s3[12][30] , \add_out_s3[12][29] ,
         \add_out_s3[12][28] , \add_out_s3[12][27] , \add_out_s3[12][26] ,
         \add_out_s3[12][25] , \add_out_s3[12][24] , \add_out_s3[12][23] ,
         \add_out_s3[12][22] , \add_out_s3[12][21] , \add_out_s3[12][20] ,
         \add_out_s3[12][19] , \add_out_s3[12][18] , \add_out_s3[12][17] ,
         \add_out_s3[12][16] , \add_out_s3[12][15] , \add_out_s3[12][14] ,
         \add_out_s3[12][13] , \add_out_s3[12][12] , \add_out_s3[12][11] ,
         \add_out_s3[12][10] , \add_out_s3[12][9] , \add_out_s3[12][8] ,
         \add_out_s3[12][7] , \add_out_s3[12][6] , \add_out_s3[12][5] ,
         \add_out_s3[12][4] , \add_out_s3[12][3] , \add_out_s3[12][2] ,
         \add_out_s3[12][1] , \add_out_s3[12][0] , \add_out_s3[11][31] ,
         \add_out_s3[11][30] , \add_out_s3[11][29] , \add_out_s3[11][28] ,
         \add_out_s3[11][27] , \add_out_s3[11][26] , \add_out_s3[11][25] ,
         \add_out_s3[11][24] , \add_out_s3[11][23] , \add_out_s3[11][22] ,
         \add_out_s3[11][21] , \add_out_s3[11][20] , \add_out_s3[11][19] ,
         \add_out_s3[11][18] , \add_out_s3[11][17] , \add_out_s3[11][16] ,
         \add_out_s3[11][15] , \add_out_s3[11][14] , \add_out_s3[11][13] ,
         \add_out_s3[11][12] , \add_out_s3[11][11] , \add_out_s3[11][10] ,
         \add_out_s3[11][9] , \add_out_s3[11][8] , \add_out_s3[11][7] ,
         \add_out_s3[11][6] , \add_out_s3[11][5] , \add_out_s3[11][4] ,
         \add_out_s3[11][3] , \add_out_s3[11][2] , \add_out_s3[11][1] ,
         \add_out_s3[11][0] , \add_out_s3[10][31] , \add_out_s3[10][30] ,
         \add_out_s3[10][29] , \add_out_s3[10][28] , \add_out_s3[10][27] ,
         \add_out_s3[10][26] , \add_out_s3[10][25] , \add_out_s3[10][24] ,
         \add_out_s3[10][23] , \add_out_s3[10][22] , \add_out_s3[10][21] ,
         \add_out_s3[10][20] , \add_out_s3[10][19] , \add_out_s3[10][18] ,
         \add_out_s3[10][17] , \add_out_s3[10][16] , \add_out_s3[10][15] ,
         \add_out_s3[10][14] , \add_out_s3[10][13] , \add_out_s3[10][12] ,
         \add_out_s3[10][11] , \add_out_s3[10][10] , \add_out_s3[10][9] ,
         \add_out_s3[10][8] , \add_out_s3[10][7] , \add_out_s3[10][6] ,
         \add_out_s3[10][5] , \add_out_s3[10][4] , \add_out_s3[10][3] ,
         \add_out_s3[10][2] , \add_out_s3[10][1] , \add_out_s3[10][0] ,
         \add_out_s3[9][31] , \add_out_s3[9][30] , \add_out_s3[9][29] ,
         \add_out_s3[9][28] , \add_out_s3[9][27] , \add_out_s3[9][26] ,
         \add_out_s3[9][25] , \add_out_s3[9][24] , \add_out_s3[9][23] ,
         \add_out_s3[9][22] , \add_out_s3[9][21] , \add_out_s3[9][20] ,
         \add_out_s3[9][19] , \add_out_s3[9][18] , \add_out_s3[9][17] ,
         \add_out_s3[9][16] , \add_out_s3[9][15] , \add_out_s3[9][14] ,
         \add_out_s3[9][13] , \add_out_s3[9][12] , \add_out_s3[9][11] ,
         \add_out_s3[9][10] , \add_out_s3[9][9] , \add_out_s3[9][8] ,
         \add_out_s3[9][7] , \add_out_s3[9][6] , \add_out_s3[9][5] ,
         \add_out_s3[9][4] , \add_out_s3[9][3] , \add_out_s3[9][2] ,
         \add_out_s3[9][1] , \add_out_s3[9][0] , \add_out_s3[8][31] ,
         \add_out_s3[8][30] , \add_out_s3[8][29] , \add_out_s3[8][28] ,
         \add_out_s3[8][27] , \add_out_s3[8][26] , \add_out_s3[8][25] ,
         \add_out_s3[8][24] , \add_out_s3[8][23] , \add_out_s3[8][22] ,
         \add_out_s3[8][21] , \add_out_s3[8][20] , \add_out_s3[8][19] ,
         \add_out_s3[8][18] , \add_out_s3[8][17] , \add_out_s3[8][16] ,
         \add_out_s3[8][15] , \add_out_s3[8][14] , \add_out_s3[8][13] ,
         \add_out_s3[8][12] , \add_out_s3[8][11] , \add_out_s3[8][10] ,
         \add_out_s3[8][9] , \add_out_s3[8][8] , \add_out_s3[8][7] ,
         \add_out_s3[8][6] , \add_out_s3[8][5] , \add_out_s3[8][4] ,
         \add_out_s3[8][3] , \add_out_s3[8][2] , \add_out_s3[8][1] ,
         \add_out_s3[8][0] , \add_out_s4[14][31] , \add_out_s4[14][30] ,
         \add_out_s4[14][29] , \add_out_s4[14][28] , \add_out_s4[14][27] ,
         \add_out_s4[14][26] , \add_out_s4[14][25] , \add_out_s4[14][24] ,
         \add_out_s4[14][23] , \add_out_s4[14][22] , \add_out_s4[14][21] ,
         \add_out_s4[14][20] , \add_out_s4[14][19] , \add_out_s4[14][18] ,
         \add_out_s4[14][17] , \add_out_s4[14][16] , \add_out_s4[14][15] ,
         \add_out_s4[14][14] , \add_out_s4[14][13] , \add_out_s4[14][12] ,
         \add_out_s4[14][11] , \add_out_s4[14][10] , \add_out_s4[14][9] ,
         \add_out_s4[14][8] , \add_out_s4[14][7] , \add_out_s4[14][6] ,
         \add_out_s4[14][5] , \add_out_s4[14][4] , \add_out_s4[14][3] ,
         \add_out_s4[14][2] , \add_out_s4[14][1] , \add_out_s4[14][0] ,
         \add_out_s4[13][31] , \add_out_s4[13][30] , \add_out_s4[13][29] ,
         \add_out_s4[13][28] , \add_out_s4[13][27] , \add_out_s4[13][26] ,
         \add_out_s4[13][25] , \add_out_s4[13][24] , \add_out_s4[13][23] ,
         \add_out_s4[13][22] , \add_out_s4[13][21] , \add_out_s4[13][20] ,
         \add_out_s4[13][19] , \add_out_s4[13][18] , \add_out_s4[13][17] ,
         \add_out_s4[13][16] , \add_out_s4[13][15] , \add_out_s4[13][14] ,
         \add_out_s4[13][13] , \add_out_s4[13][12] , \add_out_s4[13][11] ,
         \add_out_s4[13][10] , \add_out_s4[13][9] , \add_out_s4[13][8] ,
         \add_out_s4[13][7] , \add_out_s4[13][6] , \add_out_s4[13][5] ,
         \add_out_s4[13][4] , \add_out_s4[13][3] , \add_out_s4[13][2] ,
         \add_out_s4[13][1] , \add_out_s4[13][0] , \add_out_s4[12][31] ,
         \add_out_s4[12][30] , \add_out_s4[12][29] , \add_out_s4[12][28] ,
         \add_out_s4[12][27] , \add_out_s4[12][26] , \add_out_s4[12][25] ,
         \add_out_s4[12][24] , \add_out_s4[12][23] , \add_out_s4[12][22] ,
         \add_out_s4[12][21] , \add_out_s4[12][20] , \add_out_s4[12][19] ,
         \add_out_s4[12][18] , \add_out_s4[12][17] , \add_out_s4[12][16] ,
         \add_out_s4[12][15] , \add_out_s4[12][14] , \add_out_s4[12][13] ,
         \add_out_s4[12][12] , \add_out_s4[12][11] , \add_out_s4[12][10] ,
         \add_out_s4[12][9] , \add_out_s4[12][8] , \add_out_s4[12][7] ,
         \add_out_s4[12][6] , \add_out_s4[12][5] , \add_out_s4[12][4] ,
         \add_out_s4[12][3] , \add_out_s4[12][2] , \add_out_s4[12][1] ,
         \add_out_s4[12][0] , \add_out_s1[4][31] , \add_out_s1[4][30] ,
         \add_out_s1[4][29] , \add_out_s1[4][28] , \add_out_s1[4][27] ,
         \add_out_s1[4][26] , \add_out_s1[4][25] , \add_out_s1[4][24] ,
         \add_out_s1[4][23] , \add_out_s1[4][22] , \add_out_s1[4][21] ,
         \add_out_s1[4][20] , \add_out_s1[4][19] , \add_out_s1[4][18] ,
         \add_out_s1[4][17] , \add_out_s1[4][16] , \add_out_s1[4][15] ,
         \add_out_s1[4][14] , \add_out_s1[4][13] , \add_out_s1[4][12] ,
         \add_out_s1[4][11] , \add_out_s1[4][10] , \add_out_s1[4][9] ,
         \add_out_s1[4][8] , \add_out_s1[4][7] , \add_out_s1[4][6] ,
         \add_out_s1[4][5] , \add_out_s1[4][4] , \add_out_s1[4][3] ,
         \add_out_s1[4][2] , \add_out_s1[4][1] , \add_out_s1[4][0] ,
         \add_out_s1[3][31] , \add_out_s1[3][30] , \add_out_s1[3][29] ,
         \add_out_s1[3][28] , \add_out_s1[3][27] , \add_out_s1[3][26] ,
         \add_out_s1[3][25] , \add_out_s1[3][24] , \add_out_s1[3][23] ,
         \add_out_s1[3][22] , \add_out_s1[3][21] , \add_out_s1[3][20] ,
         \add_out_s1[3][19] , \add_out_s1[3][18] , \add_out_s1[3][17] ,
         \add_out_s1[3][16] , \add_out_s1[3][14] , \add_out_s1[3][13] ,
         \add_out_s1[3][12] , \add_out_s1[3][11] , \add_out_s1[3][10] ,
         \add_out_s1[3][9] , \add_out_s1[3][8] , \add_out_s1[3][7] ,
         \add_out_s1[3][6] , \add_out_s1[3][5] , \add_out_s1[3][4] ,
         \add_out_s1[3][3] , \add_out_s1[3][2] , \add_out_s1[3][1] ,
         \add_out_s1[3][0] , \add_out_s1[2][31] , \add_out_s1[2][30] ,
         \add_out_s1[2][29] , \add_out_s1[2][28] , \add_out_s1[2][27] ,
         \add_out_s1[2][26] , \add_out_s1[2][25] , \add_out_s1[2][24] ,
         \add_out_s1[2][23] , \add_out_s1[2][22] , \add_out_s1[2][21] ,
         \add_out_s1[2][20] , \add_out_s1[2][19] , \add_out_s1[2][18] ,
         \add_out_s1[2][17] , \add_out_s1[2][16] , \add_out_s1[2][15] ,
         \add_out_s1[2][14] , \add_out_s1[2][13] , \add_out_s1[2][12] ,
         \add_out_s1[2][11] , \add_out_s1[2][10] , \add_out_s1[2][9] ,
         \add_out_s1[2][8] , \add_out_s1[2][7] , \add_out_s1[2][6] ,
         \add_out_s1[2][5] , \add_out_s1[2][4] , \add_out_s1[2][3] ,
         \add_out_s1[2][2] , \add_out_s1[2][1] , \add_out_s1[2][0] ,
         \add_out_s1[1][31] , \add_out_s1[1][30] , \add_out_s1[1][29] ,
         \add_out_s1[1][28] , \add_out_s1[1][27] , \add_out_s1[1][26] ,
         \add_out_s1[1][25] , \add_out_s1[1][23] , \add_out_s1[1][22] ,
         \add_out_s1[1][21] , \add_out_s1[1][20] , \add_out_s1[1][19] ,
         \add_out_s1[1][18] , \add_out_s1[1][17] , \add_out_s1[1][16] ,
         \add_out_s1[1][15] , \add_out_s1[1][14] , \add_out_s1[1][13] ,
         \add_out_s1[1][12] , \add_out_s1[1][11] , \add_out_s1[1][10] ,
         \add_out_s1[1][9] , \add_out_s1[1][8] , \add_out_s1[1][7] ,
         \add_out_s1[1][6] , \add_out_s1[1][5] , \add_out_s1[1][4] ,
         \add_out_s1[1][3] , \add_out_s1[1][2] , \add_out_s1[1][1] ,
         \add_out_s1[1][0] , \add_out_s1[0][31] , \add_out_s1[0][30] ,
         \add_out_s1[0][29] , \add_out_s1[0][28] , \add_out_s1[0][27] ,
         \add_out_s1[0][26] , \add_out_s1[0][25] , \add_out_s1[0][24] ,
         \add_out_s1[0][23] , \add_out_s1[0][22] , \add_out_s1[0][21] ,
         \add_out_s1[0][20] , \add_out_s1[0][19] , \add_out_s1[0][18] ,
         \add_out_s1[0][17] , \add_out_s1[0][16] , \add_out_s1[0][15] ,
         \add_out_s1[0][14] , \add_out_s1[0][13] , \add_out_s1[0][12] ,
         \add_out_s1[0][11] , \add_out_s1[0][10] , \add_out_s1[0][9] ,
         \add_out_s1[0][8] , \add_out_s1[0][7] , \add_out_s1[0][6] ,
         \add_out_s1[0][5] , \add_out_s1[0][4] , \add_out_s1[0][3] ,
         \add_out_s1[0][2] , \add_out_s1[0][1] , \add_out_s1[0][0] ,
         \add_out_s2[8][31] , \add_out_s2[8][30] , \add_out_s2[8][29] ,
         \add_out_s2[8][28] , \add_out_s2[8][27] , \add_out_s2[8][26] ,
         \add_out_s2[8][25] , \add_out_s2[8][24] , \add_out_s2[8][23] ,
         \add_out_s2[8][22] , \add_out_s2[8][21] , \add_out_s2[8][20] ,
         \add_out_s2[8][19] , \add_out_s2[8][18] , \add_out_s2[8][17] ,
         \add_out_s2[8][16] , \add_out_s2[8][15] , \add_out_s2[8][14] ,
         \add_out_s2[8][13] , \add_out_s2[8][12] , \add_out_s2[8][11] ,
         \add_out_s2[8][10] , \add_out_s2[8][9] , \add_out_s2[8][8] ,
         \add_out_s2[8][7] , \add_out_s2[8][6] , \add_out_s2[8][5] ,
         \add_out_s2[8][4] , \add_out_s2[8][3] , \add_out_s2[8][2] ,
         \add_out_s2[8][1] , \add_out_s2[8][0] , \A_shifted[-32][62] ,
         \A_shifted[-32][61] , \A_shifted[-32][60] , \A_shifted[-32][59] ,
         \A_shifted[-32][58] , \A_shifted[-32][57] , \A_shifted[-32][56] ,
         \A_shifted[-32][55] , \A_shifted[-32][54] , \A_shifted[-32][53] ,
         \A_shifted[-32][52] , \A_shifted[-32][51] , \A_shifted[-32][50] ,
         \A_shifted[-32][49] , \A_shifted[-32][48] , \A_shifted[-32][47] ,
         \A_shifted[-32][46] , \A_shifted[-32][45] , \A_shifted[-32][44] ,
         \A_shifted[-32][43] , \A_shifted[-32][42] , \A_shifted[-32][41] ,
         \A_shifted[-32][40] , \A_shifted[-32][39] , \A_shifted[-32][38] ,
         \A_shifted[-32][37] , \A_shifted[-32][36] , \A_shifted[-32][35] ,
         \A_shifted[-32][34] , \A_shifted[-32][33] , \A_shifted[-32][32] ,
         \mux_out[7][31] , \mux_out[7][30] , \mux_out[7][29] ,
         \mux_out[7][28] , \mux_out[7][27] , \mux_out[7][26] ,
         \mux_out[7][25] , \mux_out[7][24] , \mux_out[7][23] ,
         \mux_out[7][22] , \mux_out[7][21] , \mux_out[7][20] ,
         \mux_out[7][19] , \mux_out[7][18] , \mux_out[7][17] ,
         \mux_out[7][16] , \mux_out[7][15] , \mux_out[7][14] ,
         \mux_out[6][31] , \mux_out[6][30] , \mux_out[6][29] ,
         \mux_out[6][28] , \mux_out[6][27] , \mux_out[6][26] ,
         \mux_out[6][25] , \mux_out[6][24] , \mux_out[6][23] ,
         \mux_out[6][22] , \mux_out[6][21] , \mux_out[6][20] ,
         \mux_out[6][19] , \mux_out[6][18] , \mux_out[6][17] ,
         \mux_out[6][16] , \mux_out[6][15] , \mux_out[6][14] ,
         \mux_out[6][13] , \mux_out[6][12] , \mux_out[5][31] ,
         \mux_out[5][30] , \mux_out[5][29] , \mux_out[5][28] ,
         \mux_out[5][27] , \mux_out[5][26] , \mux_out[5][25] ,
         \mux_out[5][24] , \mux_out[5][23] , \mux_out[5][22] ,
         \mux_out[5][21] , \mux_out[5][19] , \mux_out[5][18] ,
         \mux_out[5][17] , \mux_out[5][16] , \mux_out[5][15] ,
         \mux_out[5][14] , \mux_out[5][13] , \mux_out[5][12] ,
         \mux_out[5][11] , \mux_out[5][10] , \mux_out[4][31] ,
         \mux_out[4][30] , \mux_out[4][29] , \mux_out[4][28] ,
         \mux_out[4][27] , \mux_out[4][26] , \mux_out[4][25] ,
         \mux_out[4][24] , \mux_out[4][23] , \mux_out[4][22] ,
         \mux_out[4][21] , \mux_out[4][20] , \mux_out[4][19] ,
         \mux_out[4][18] , \mux_out[4][17] , \mux_out[4][16] ,
         \mux_out[4][15] , \mux_out[4][14] , \mux_out[4][13] ,
         \mux_out[4][12] , \mux_out[4][11] , \mux_out[4][10] , \mux_out[4][9] ,
         \mux_out[4][8] , \mux_out[3][31] , \mux_out[3][30] , \mux_out[3][29] ,
         \mux_out[3][28] , \mux_out[3][27] , \mux_out[3][26] ,
         \mux_out[3][25] , \mux_out[3][24] , \mux_out[3][23] ,
         \mux_out[3][22] , \mux_out[3][21] , \mux_out[3][20] ,
         \mux_out[3][19] , \mux_out[3][18] , \mux_out[3][17] ,
         \mux_out[3][16] , \mux_out[3][15] , \mux_out[3][14] ,
         \mux_out[3][13] , \mux_out[3][12] , \mux_out[3][11] ,
         \mux_out[3][10] , \mux_out[3][9] , \mux_out[3][8] , \mux_out[3][7] ,
         \mux_out[3][6] , \mux_out[2][31] , \mux_out[2][30] , \mux_out[2][29] ,
         \mux_out[2][28] , \mux_out[2][27] , \mux_out[2][26] ,
         \mux_out[2][25] , \mux_out[2][24] , \mux_out[2][23] ,
         \mux_out[2][22] , \mux_out[2][21] , \mux_out[2][20] ,
         \mux_out[2][19] , \mux_out[2][18] , \mux_out[2][17] ,
         \mux_out[2][16] , \mux_out[2][15] , \mux_out[2][14] ,
         \mux_out[2][13] , \mux_out[2][12] , \mux_out[2][11] ,
         \mux_out[2][10] , \mux_out[2][9] , \mux_out[2][8] , \mux_out[2][7] ,
         \mux_out[2][6] , \mux_out[2][5] , \mux_out[2][4] , \mux_out[1][31] ,
         \mux_out[1][30] , \mux_out[1][29] , \mux_out[1][28] ,
         \mux_out[1][27] , \mux_out[1][26] , \mux_out[1][25] ,
         \mux_out[1][24] , \mux_out[1][23] , \mux_out[1][22] ,
         \mux_out[1][21] , \mux_out[1][20] , \mux_out[1][19] ,
         \mux_out[1][18] , \mux_out[1][17] , \mux_out[1][16] ,
         \mux_out[1][15] , \mux_out[1][14] , \mux_out[1][13] ,
         \mux_out[1][12] , \mux_out[1][11] , \mux_out[1][10] , \mux_out[1][9] ,
         \mux_out[1][8] , \mux_out[1][7] , \mux_out[1][6] , \mux_out[1][5] ,
         \mux_out[1][4] , \mux_out[1][3] , \mux_out[1][2] , \mux_out[15][31] ,
         \mux_out[15][30] , \mux_out[14][31] , \mux_out[14][30] ,
         \mux_out[14][29] , \mux_out[14][28] , \mux_out[13][31] ,
         \mux_out[13][30] , \mux_out[13][29] , \mux_out[13][28] ,
         \mux_out[13][27] , \mux_out[13][26] , \mux_out[12][31] ,
         \mux_out[12][30] , \mux_out[12][29] , \mux_out[12][28] ,
         \mux_out[12][27] , \mux_out[12][26] , \mux_out[12][25] ,
         \mux_out[12][24] , \mux_out[11][31] , \mux_out[11][30] ,
         \mux_out[11][29] , \mux_out[11][28] , \mux_out[11][27] ,
         \mux_out[11][26] , \mux_out[11][25] , \mux_out[11][24] ,
         \mux_out[11][23] , \mux_out[11][22] , \mux_out[10][31] ,
         \mux_out[10][30] , \mux_out[10][29] , \mux_out[10][28] ,
         \mux_out[10][27] , \mux_out[10][26] , \mux_out[10][25] ,
         \mux_out[10][24] , \mux_out[10][23] , \mux_out[10][22] ,
         \mux_out[10][21] , \mux_out[10][20] , \mux_out[9][31] ,
         \mux_out[9][30] , \mux_out[9][29] , \mux_out[9][28] ,
         \mux_out[9][27] , \mux_out[9][26] , \mux_out[9][25] ,
         \mux_out[9][24] , \mux_out[9][23] , \mux_out[9][22] ,
         \mux_out[9][21] , \mux_out[9][20] , \mux_out[9][19] ,
         \mux_out[9][18] , \mux_out[8][31] , \mux_out[8][30] ,
         \mux_out[8][29] , \mux_out[8][28] , \mux_out[8][27] ,
         \mux_out[8][26] , \mux_out[8][25] , \mux_out[8][24] ,
         \mux_out[8][23] , \mux_out[8][22] , \mux_out[8][21] ,
         \mux_out[8][20] , \mux_out[8][19] , \mux_out[8][18] ,
         \mux_out[8][17] , \mux_out[8][16] , \encoder_out[15][2] ,
         \encoder_out[15][1] , \encoder_out[15][0] , \encoder_out[14][2] ,
         \encoder_out[14][1] , \encoder_out[14][0] , \encoder_out[13][2] ,
         \encoder_out[13][1] , \encoder_out[13][0] , \encoder_out[12][2] ,
         \encoder_out[12][1] , \encoder_out[12][0] , \encoder_out[11][2] ,
         \encoder_out[11][1] , \encoder_out[11][0] , \encoder_out[10][2] ,
         \encoder_out[10][1] , \encoder_out[10][0] , \encoder_out[9][2] ,
         \encoder_out[9][1] , \encoder_out[9][0] , \encoder_out[8][2] ,
         \encoder_out[8][1] , \encoder_out[8][0] , \encoder_out[7][2] ,
         \encoder_out[7][1] , \encoder_out[7][0] , \encoder_out[6][2] ,
         \encoder_out[6][1] , \encoder_out[6][0] , \encoder_out[5][2] ,
         \encoder_out[5][1] , \encoder_out[5][0] , \encoder_out[4][2] ,
         \encoder_out[4][1] , \encoder_out[4][0] , \encoder_out[3][2] ,
         \encoder_out[3][1] , \encoder_out[3][0] , \encoder_out[2][2] ,
         \encoder_out[2][1] , \encoder_out[2][0] , \encoder_out[1][2] ,
         \encoder_out[1][1] , \encoder_out[1][0] , \encoder_out[0][2] ,
         \encoder_out[0][1] , \encoder_out[0][0] , net18822, net18832,
         net18842, \sub_x_1/B[23] , \sub_x_1/B[22] , \sub_x_1/B[21] ,
         \sub_x_1/B[17] , \sub_x_1/B[15] , \sub_x_1/n29 , \sub_x_1/n26 ,
         \sub_x_1/n25 , \sub_x_1/n24 , \sub_x_1/n21 , \sub_x_1/n19 ,
         \sub_x_1/n17 , \sub_x_1/n16 , \sub_x_1/n15 , \sub_x_1/n11 ,
         \sub_x_1/n10 , \sub_x_1/n9 , \sub_x_1/n8 , \sub_x_1/n7 , \sub_x_1/n6 ,
         \sub_x_1/n5 , \sub_x_1/n4 , \sub_x_1/n3 , \sub_x_1/n2 , n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n12, n13, n14, n15, n16, n17, n18, n19, n22,
         n23, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106, SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        SYNOPSYS_UNCONNECTED__118, SYNOPSYS_UNCONNECTED__119, 
        SYNOPSYS_UNCONNECTED__120, SYNOPSYS_UNCONNECTED__121, 
        SYNOPSYS_UNCONNECTED__122, SYNOPSYS_UNCONNECTED__123, 
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        SYNOPSYS_UNCONNECTED__126, SYNOPSYS_UNCONNECTED__127, 
        SYNOPSYS_UNCONNECTED__128, SYNOPSYS_UNCONNECTED__129, 
        SYNOPSYS_UNCONNECTED__130, SYNOPSYS_UNCONNECTED__131, 
        SYNOPSYS_UNCONNECTED__132, SYNOPSYS_UNCONNECTED__133, 
        SYNOPSYS_UNCONNECTED__134, SYNOPSYS_UNCONNECTED__135, 
        SYNOPSYS_UNCONNECTED__136, SYNOPSYS_UNCONNECTED__137, 
        SYNOPSYS_UNCONNECTED__138, SYNOPSYS_UNCONNECTED__139, 
        SYNOPSYS_UNCONNECTED__140, SYNOPSYS_UNCONNECTED__141, 
        SYNOPSYS_UNCONNECTED__142, SYNOPSYS_UNCONNECTED__143, 
        SYNOPSYS_UNCONNECTED__144, SYNOPSYS_UNCONNECTED__145, 
        SYNOPSYS_UNCONNECTED__146, SYNOPSYS_UNCONNECTED__147, 
        SYNOPSYS_UNCONNECTED__148, SYNOPSYS_UNCONNECTED__149, 
        SYNOPSYS_UNCONNECTED__150, SYNOPSYS_UNCONNECTED__151, 
        SYNOPSYS_UNCONNECTED__152, SYNOPSYS_UNCONNECTED__153, 
        SYNOPSYS_UNCONNECTED__154, SYNOPSYS_UNCONNECTED__155, 
        SYNOPSYS_UNCONNECTED__156, SYNOPSYS_UNCONNECTED__157, 
        SYNOPSYS_UNCONNECTED__158, SYNOPSYS_UNCONNECTED__159, 
        SYNOPSYS_UNCONNECTED__160, SYNOPSYS_UNCONNECTED__161, 
        SYNOPSYS_UNCONNECTED__162, SYNOPSYS_UNCONNECTED__163, 
        SYNOPSYS_UNCONNECTED__164, SYNOPSYS_UNCONNECTED__165, 
        SYNOPSYS_UNCONNECTED__166, SYNOPSYS_UNCONNECTED__167, 
        SYNOPSYS_UNCONNECTED__168, SYNOPSYS_UNCONNECTED__169, 
        SYNOPSYS_UNCONNECTED__170, SYNOPSYS_UNCONNECTED__171, 
        SYNOPSYS_UNCONNECTED__172, SYNOPSYS_UNCONNECTED__173, 
        SYNOPSYS_UNCONNECTED__174, SYNOPSYS_UNCONNECTED__175, 
        SYNOPSYS_UNCONNECTED__176, SYNOPSYS_UNCONNECTED__177, 
        SYNOPSYS_UNCONNECTED__178, SYNOPSYS_UNCONNECTED__179, 
        SYNOPSYS_UNCONNECTED__180, SYNOPSYS_UNCONNECTED__181, 
        SYNOPSYS_UNCONNECTED__182, SYNOPSYS_UNCONNECTED__183, 
        SYNOPSYS_UNCONNECTED__184, SYNOPSYS_UNCONNECTED__185, 
        SYNOPSYS_UNCONNECTED__186, SYNOPSYS_UNCONNECTED__187, 
        SYNOPSYS_UNCONNECTED__188, SYNOPSYS_UNCONNECTED__189, 
        SYNOPSYS_UNCONNECTED__190, SYNOPSYS_UNCONNECTED__191, 
        SYNOPSYS_UNCONNECTED__192, SYNOPSYS_UNCONNECTED__193, 
        SYNOPSYS_UNCONNECTED__194, SYNOPSYS_UNCONNECTED__195, 
        SYNOPSYS_UNCONNECTED__196, SYNOPSYS_UNCONNECTED__197, 
        SYNOPSYS_UNCONNECTED__198, SYNOPSYS_UNCONNECTED__199, 
        SYNOPSYS_UNCONNECTED__200, SYNOPSYS_UNCONNECTED__201, 
        SYNOPSYS_UNCONNECTED__202, SYNOPSYS_UNCONNECTED__203, 
        SYNOPSYS_UNCONNECTED__204, SYNOPSYS_UNCONNECTED__205, 
        SYNOPSYS_UNCONNECTED__206, SYNOPSYS_UNCONNECTED__207, 
        SYNOPSYS_UNCONNECTED__208, SYNOPSYS_UNCONNECTED__209, 
        SYNOPSYS_UNCONNECTED__210, SYNOPSYS_UNCONNECTED__211, 
        SYNOPSYS_UNCONNECTED__212, SYNOPSYS_UNCONNECTED__213, 
        SYNOPSYS_UNCONNECTED__214, SYNOPSYS_UNCONNECTED__215, 
        SYNOPSYS_UNCONNECTED__216, SYNOPSYS_UNCONNECTED__217, 
        SYNOPSYS_UNCONNECTED__218, SYNOPSYS_UNCONNECTED__219, 
        SYNOPSYS_UNCONNECTED__220, SYNOPSYS_UNCONNECTED__221, 
        SYNOPSYS_UNCONNECTED__222, SYNOPSYS_UNCONNECTED__223, 
        SYNOPSYS_UNCONNECTED__224, SYNOPSYS_UNCONNECTED__225, 
        SYNOPSYS_UNCONNECTED__226, SYNOPSYS_UNCONNECTED__227, 
        SYNOPSYS_UNCONNECTED__228, SYNOPSYS_UNCONNECTED__229, 
        SYNOPSYS_UNCONNECTED__230, SYNOPSYS_UNCONNECTED__231, 
        SYNOPSYS_UNCONNECTED__232, SYNOPSYS_UNCONNECTED__233, 
        SYNOPSYS_UNCONNECTED__234, SYNOPSYS_UNCONNECTED__235, 
        SYNOPSYS_UNCONNECTED__236, SYNOPSYS_UNCONNECTED__237, 
        SYNOPSYS_UNCONNECTED__238, SYNOPSYS_UNCONNECTED__239, 
        SYNOPSYS_UNCONNECTED__240, SYNOPSYS_UNCONNECTED__241, 
        SYNOPSYS_UNCONNECTED__242, SYNOPSYS_UNCONNECTED__243, 
        SYNOPSYS_UNCONNECTED__244, SYNOPSYS_UNCONNECTED__245, 
        SYNOPSYS_UNCONNECTED__246, SYNOPSYS_UNCONNECTED__247, 
        SYNOPSYS_UNCONNECTED__248, SYNOPSYS_UNCONNECTED__249, 
        SYNOPSYS_UNCONNECTED__250, SYNOPSYS_UNCONNECTED__251, 
        SYNOPSYS_UNCONNECTED__252, SYNOPSYS_UNCONNECTED__253, 
        SYNOPSYS_UNCONNECTED__254, SYNOPSYS_UNCONNECTED__255, 
        SYNOPSYS_UNCONNECTED__256, SYNOPSYS_UNCONNECTED__257, 
        SYNOPSYS_UNCONNECTED__258, SYNOPSYS_UNCONNECTED__259, 
        SYNOPSYS_UNCONNECTED__260, SYNOPSYS_UNCONNECTED__261, 
        SYNOPSYS_UNCONNECTED__262, SYNOPSYS_UNCONNECTED__263, 
        SYNOPSYS_UNCONNECTED__264, SYNOPSYS_UNCONNECTED__265, 
        SYNOPSYS_UNCONNECTED__266, SYNOPSYS_UNCONNECTED__267, 
        SYNOPSYS_UNCONNECTED__268, SYNOPSYS_UNCONNECTED__269, 
        SYNOPSYS_UNCONNECTED__270, SYNOPSYS_UNCONNECTED__271, 
        SYNOPSYS_UNCONNECTED__272, SYNOPSYS_UNCONNECTED__273, 
        SYNOPSYS_UNCONNECTED__274, SYNOPSYS_UNCONNECTED__275, 
        SYNOPSYS_UNCONNECTED__276, SYNOPSYS_UNCONNECTED__277, 
        SYNOPSYS_UNCONNECTED__278, SYNOPSYS_UNCONNECTED__279, 
        SYNOPSYS_UNCONNECTED__280, SYNOPSYS_UNCONNECTED__281, 
        SYNOPSYS_UNCONNECTED__282, SYNOPSYS_UNCONNECTED__283, 
        SYNOPSYS_UNCONNECTED__284, SYNOPSYS_UNCONNECTED__285, 
        SYNOPSYS_UNCONNECTED__286, SYNOPSYS_UNCONNECTED__287, 
        SYNOPSYS_UNCONNECTED__288, SYNOPSYS_UNCONNECTED__289, 
        SYNOPSYS_UNCONNECTED__290, SYNOPSYS_UNCONNECTED__291, 
        SYNOPSYS_UNCONNECTED__292, SYNOPSYS_UNCONNECTED__293, 
        SYNOPSYS_UNCONNECTED__294, SYNOPSYS_UNCONNECTED__295, 
        SYNOPSYS_UNCONNECTED__296, SYNOPSYS_UNCONNECTED__297, 
        SYNOPSYS_UNCONNECTED__298, SYNOPSYS_UNCONNECTED__299, 
        SYNOPSYS_UNCONNECTED__300, SYNOPSYS_UNCONNECTED__301, 
        SYNOPSYS_UNCONNECTED__302, SYNOPSYS_UNCONNECTED__303, 
        SYNOPSYS_UNCONNECTED__304, SYNOPSYS_UNCONNECTED__305, 
        SYNOPSYS_UNCONNECTED__306, SYNOPSYS_UNCONNECTED__307, 
        SYNOPSYS_UNCONNECTED__308, SYNOPSYS_UNCONNECTED__309, 
        SYNOPSYS_UNCONNECTED__310, SYNOPSYS_UNCONNECTED__311, 
        SYNOPSYS_UNCONNECTED__312, SYNOPSYS_UNCONNECTED__313, 
        SYNOPSYS_UNCONNECTED__314, SYNOPSYS_UNCONNECTED__315, 
        SYNOPSYS_UNCONNECTED__316, SYNOPSYS_UNCONNECTED__317, 
        SYNOPSYS_UNCONNECTED__318, SYNOPSYS_UNCONNECTED__319, 
        SYNOPSYS_UNCONNECTED__320, SYNOPSYS_UNCONNECTED__321, 
        SYNOPSYS_UNCONNECTED__322, SYNOPSYS_UNCONNECTED__323, 
        SYNOPSYS_UNCONNECTED__324, SYNOPSYS_UNCONNECTED__325, 
        SYNOPSYS_UNCONNECTED__326, SYNOPSYS_UNCONNECTED__327, 
        SYNOPSYS_UNCONNECTED__328, SYNOPSYS_UNCONNECTED__329, 
        SYNOPSYS_UNCONNECTED__330, SYNOPSYS_UNCONNECTED__331, 
        SYNOPSYS_UNCONNECTED__332, SYNOPSYS_UNCONNECTED__333, 
        SYNOPSYS_UNCONNECTED__334, SYNOPSYS_UNCONNECTED__335, 
        SYNOPSYS_UNCONNECTED__336, SYNOPSYS_UNCONNECTED__337, 
        SYNOPSYS_UNCONNECTED__338, SYNOPSYS_UNCONNECTED__339, 
        SYNOPSYS_UNCONNECTED__340, SYNOPSYS_UNCONNECTED__341, 
        SYNOPSYS_UNCONNECTED__342, SYNOPSYS_UNCONNECTED__343, 
        SYNOPSYS_UNCONNECTED__344, SYNOPSYS_UNCONNECTED__345, 
        SYNOPSYS_UNCONNECTED__346, SYNOPSYS_UNCONNECTED__347, 
        SYNOPSYS_UNCONNECTED__348, SYNOPSYS_UNCONNECTED__349, 
        SYNOPSYS_UNCONNECTED__350, SYNOPSYS_UNCONNECTED__351, 
        SYNOPSYS_UNCONNECTED__352, SYNOPSYS_UNCONNECTED__353, 
        SYNOPSYS_UNCONNECTED__354, SYNOPSYS_UNCONNECTED__355, 
        SYNOPSYS_UNCONNECTED__356, SYNOPSYS_UNCONNECTED__357, 
        SYNOPSYS_UNCONNECTED__358, SYNOPSYS_UNCONNECTED__359, 
        SYNOPSYS_UNCONNECTED__360, SYNOPSYS_UNCONNECTED__361, 
        SYNOPSYS_UNCONNECTED__362, SYNOPSYS_UNCONNECTED__363, 
        SYNOPSYS_UNCONNECTED__364, SYNOPSYS_UNCONNECTED__365, 
        SYNOPSYS_UNCONNECTED__366, SYNOPSYS_UNCONNECTED__367, 
        SYNOPSYS_UNCONNECTED__368, SYNOPSYS_UNCONNECTED__369, 
        SYNOPSYS_UNCONNECTED__370, SYNOPSYS_UNCONNECTED__371, 
        SYNOPSYS_UNCONNECTED__372, SYNOPSYS_UNCONNECTED__373, 
        SYNOPSYS_UNCONNECTED__374, SYNOPSYS_UNCONNECTED__375, 
        SYNOPSYS_UNCONNECTED__376, SYNOPSYS_UNCONNECTED__377, 
        SYNOPSYS_UNCONNECTED__378, SYNOPSYS_UNCONNECTED__379, 
        SYNOPSYS_UNCONNECTED__380, SYNOPSYS_UNCONNECTED__381, 
        SYNOPSYS_UNCONNECTED__382, SYNOPSYS_UNCONNECTED__383, 
        SYNOPSYS_UNCONNECTED__384, SYNOPSYS_UNCONNECTED__385, 
        SYNOPSYS_UNCONNECTED__386, SYNOPSYS_UNCONNECTED__387, 
        SYNOPSYS_UNCONNECTED__388, SYNOPSYS_UNCONNECTED__389, 
        SYNOPSYS_UNCONNECTED__390, SYNOPSYS_UNCONNECTED__391, 
        SYNOPSYS_UNCONNECTED__392, SYNOPSYS_UNCONNECTED__393, 
        SYNOPSYS_UNCONNECTED__394, SYNOPSYS_UNCONNECTED__395, 
        SYNOPSYS_UNCONNECTED__396, SYNOPSYS_UNCONNECTED__397, 
        SYNOPSYS_UNCONNECTED__398, SYNOPSYS_UNCONNECTED__399, 
        SYNOPSYS_UNCONNECTED__400, SYNOPSYS_UNCONNECTED__401, 
        SYNOPSYS_UNCONNECTED__402, SYNOPSYS_UNCONNECTED__403, 
        SYNOPSYS_UNCONNECTED__404, SYNOPSYS_UNCONNECTED__405, 
        SYNOPSYS_UNCONNECTED__406, SYNOPSYS_UNCONNECTED__407, 
        SYNOPSYS_UNCONNECTED__408, SYNOPSYS_UNCONNECTED__409, 
        SYNOPSYS_UNCONNECTED__410, SYNOPSYS_UNCONNECTED__411, 
        SYNOPSYS_UNCONNECTED__412, SYNOPSYS_UNCONNECTED__413, 
        SYNOPSYS_UNCONNECTED__414, SYNOPSYS_UNCONNECTED__415, 
        SYNOPSYS_UNCONNECTED__416, SYNOPSYS_UNCONNECTED__417, 
        SYNOPSYS_UNCONNECTED__418, SYNOPSYS_UNCONNECTED__419, 
        SYNOPSYS_UNCONNECTED__420, SYNOPSYS_UNCONNECTED__421, 
        SYNOPSYS_UNCONNECTED__422, SYNOPSYS_UNCONNECTED__423, 
        SYNOPSYS_UNCONNECTED__424, SYNOPSYS_UNCONNECTED__425, 
        SYNOPSYS_UNCONNECTED__426, SYNOPSYS_UNCONNECTED__427, 
        SYNOPSYS_UNCONNECTED__428, SYNOPSYS_UNCONNECTED__429, 
        SYNOPSYS_UNCONNECTED__430, SYNOPSYS_UNCONNECTED__431, 
        SYNOPSYS_UNCONNECTED__432, SYNOPSYS_UNCONNECTED__433, 
        SYNOPSYS_UNCONNECTED__434, SYNOPSYS_UNCONNECTED__435, 
        SYNOPSYS_UNCONNECTED__436, SYNOPSYS_UNCONNECTED__437, 
        SYNOPSYS_UNCONNECTED__438, SYNOPSYS_UNCONNECTED__439, 
        SYNOPSYS_UNCONNECTED__440, SYNOPSYS_UNCONNECTED__441, 
        SYNOPSYS_UNCONNECTED__442, SYNOPSYS_UNCONNECTED__443, 
        SYNOPSYS_UNCONNECTED__444, SYNOPSYS_UNCONNECTED__445, 
        SYNOPSYS_UNCONNECTED__446, SYNOPSYS_UNCONNECTED__447, 
        SYNOPSYS_UNCONNECTED__448, SYNOPSYS_UNCONNECTED__449, 
        SYNOPSYS_UNCONNECTED__450, SYNOPSYS_UNCONNECTED__451, 
        SYNOPSYS_UNCONNECTED__452, SYNOPSYS_UNCONNECTED__453, 
        SYNOPSYS_UNCONNECTED__454, SYNOPSYS_UNCONNECTED__455, 
        SYNOPSYS_UNCONNECTED__456, SYNOPSYS_UNCONNECTED__457, 
        SYNOPSYS_UNCONNECTED__458, SYNOPSYS_UNCONNECTED__459, 
        SYNOPSYS_UNCONNECTED__460, SYNOPSYS_UNCONNECTED__461, 
        SYNOPSYS_UNCONNECTED__462, SYNOPSYS_UNCONNECTED__463, 
        SYNOPSYS_UNCONNECTED__464, SYNOPSYS_UNCONNECTED__465, 
        SYNOPSYS_UNCONNECTED__466, SYNOPSYS_UNCONNECTED__467, 
        SYNOPSYS_UNCONNECTED__468, SYNOPSYS_UNCONNECTED__469, 
        SYNOPSYS_UNCONNECTED__470, SYNOPSYS_UNCONNECTED__471, 
        SYNOPSYS_UNCONNECTED__472, SYNOPSYS_UNCONNECTED__473, 
        SYNOPSYS_UNCONNECTED__474, SYNOPSYS_UNCONNECTED__475, 
        SYNOPSYS_UNCONNECTED__476, SYNOPSYS_UNCONNECTED__477, 
        SYNOPSYS_UNCONNECTED__478, SYNOPSYS_UNCONNECTED__479, 
        SYNOPSYS_UNCONNECTED__480, SYNOPSYS_UNCONNECTED__481, 
        SYNOPSYS_UNCONNECTED__482, SYNOPSYS_UNCONNECTED__483, 
        SYNOPSYS_UNCONNECTED__484, SYNOPSYS_UNCONNECTED__485, 
        SYNOPSYS_UNCONNECTED__486, SYNOPSYS_UNCONNECTED__487, 
        SYNOPSYS_UNCONNECTED__488, SYNOPSYS_UNCONNECTED__489, 
        SYNOPSYS_UNCONNECTED__490, SYNOPSYS_UNCONNECTED__491, 
        SYNOPSYS_UNCONNECTED__492, SYNOPSYS_UNCONNECTED__493, 
        SYNOPSYS_UNCONNECTED__494, SYNOPSYS_UNCONNECTED__495, 
        SYNOPSYS_UNCONNECTED__496, SYNOPSYS_UNCONNECTED__497, 
        SYNOPSYS_UNCONNECTED__498, SYNOPSYS_UNCONNECTED__499, 
        SYNOPSYS_UNCONNECTED__500, SYNOPSYS_UNCONNECTED__501, 
        SYNOPSYS_UNCONNECTED__502, SYNOPSYS_UNCONNECTED__503, 
        SYNOPSYS_UNCONNECTED__504, SYNOPSYS_UNCONNECTED__505, 
        SYNOPSYS_UNCONNECTED__506, SYNOPSYS_UNCONNECTED__507, 
        SYNOPSYS_UNCONNECTED__508, SYNOPSYS_UNCONNECTED__509, 
        SYNOPSYS_UNCONNECTED__510, SYNOPSYS_UNCONNECTED__511, 
        SYNOPSYS_UNCONNECTED__512, SYNOPSYS_UNCONNECTED__513, 
        SYNOPSYS_UNCONNECTED__514, SYNOPSYS_UNCONNECTED__515, 
        SYNOPSYS_UNCONNECTED__516, SYNOPSYS_UNCONNECTED__517, 
        SYNOPSYS_UNCONNECTED__518, SYNOPSYS_UNCONNECTED__519, 
        SYNOPSYS_UNCONNECTED__520, SYNOPSYS_UNCONNECTED__521, 
        SYNOPSYS_UNCONNECTED__522, SYNOPSYS_UNCONNECTED__523, 
        SYNOPSYS_UNCONNECTED__524, SYNOPSYS_UNCONNECTED__525, 
        SYNOPSYS_UNCONNECTED__526, SYNOPSYS_UNCONNECTED__527, 
        SYNOPSYS_UNCONNECTED__528, SYNOPSYS_UNCONNECTED__529, 
        SYNOPSYS_UNCONNECTED__530, SYNOPSYS_UNCONNECTED__531, 
        SYNOPSYS_UNCONNECTED__532, SYNOPSYS_UNCONNECTED__533, 
        SYNOPSYS_UNCONNECTED__534, SYNOPSYS_UNCONNECTED__535, 
        SYNOPSYS_UNCONNECTED__536, SYNOPSYS_UNCONNECTED__537, 
        SYNOPSYS_UNCONNECTED__538, SYNOPSYS_UNCONNECTED__539, 
        SYNOPSYS_UNCONNECTED__540, SYNOPSYS_UNCONNECTED__541, 
        SYNOPSYS_UNCONNECTED__542, SYNOPSYS_UNCONNECTED__543, 
        SYNOPSYS_UNCONNECTED__544, SYNOPSYS_UNCONNECTED__545, 
        SYNOPSYS_UNCONNECTED__546, SYNOPSYS_UNCONNECTED__547, 
        SYNOPSYS_UNCONNECTED__548, SYNOPSYS_UNCONNECTED__549, 
        SYNOPSYS_UNCONNECTED__550, SYNOPSYS_UNCONNECTED__551, 
        SYNOPSYS_UNCONNECTED__552, SYNOPSYS_UNCONNECTED__553, 
        SYNOPSYS_UNCONNECTED__554, SYNOPSYS_UNCONNECTED__555, 
        SYNOPSYS_UNCONNECTED__556, SYNOPSYS_UNCONNECTED__557, 
        SYNOPSYS_UNCONNECTED__558, SYNOPSYS_UNCONNECTED__559, 
        SYNOPSYS_UNCONNECTED__560, SYNOPSYS_UNCONNECTED__561, 
        SYNOPSYS_UNCONNECTED__562, SYNOPSYS_UNCONNECTED__563, 
        SYNOPSYS_UNCONNECTED__564, SYNOPSYS_UNCONNECTED__565, 
        SYNOPSYS_UNCONNECTED__566, SYNOPSYS_UNCONNECTED__567, 
        SYNOPSYS_UNCONNECTED__568, SYNOPSYS_UNCONNECTED__569, 
        SYNOPSYS_UNCONNECTED__570, SYNOPSYS_UNCONNECTED__571, 
        SYNOPSYS_UNCONNECTED__572, SYNOPSYS_UNCONNECTED__573, 
        SYNOPSYS_UNCONNECTED__574, SYNOPSYS_UNCONNECTED__575, 
        SYNOPSYS_UNCONNECTED__576, SYNOPSYS_UNCONNECTED__577, 
        SYNOPSYS_UNCONNECTED__578, SYNOPSYS_UNCONNECTED__579, 
        SYNOPSYS_UNCONNECTED__580, SYNOPSYS_UNCONNECTED__581, 
        SYNOPSYS_UNCONNECTED__582, SYNOPSYS_UNCONNECTED__583, 
        SYNOPSYS_UNCONNECTED__584, SYNOPSYS_UNCONNECTED__585, 
        SYNOPSYS_UNCONNECTED__586, SYNOPSYS_UNCONNECTED__587, 
        SYNOPSYS_UNCONNECTED__588, SYNOPSYS_UNCONNECTED__589, 
        SYNOPSYS_UNCONNECTED__590, SYNOPSYS_UNCONNECTED__591, 
        SYNOPSYS_UNCONNECTED__592, SYNOPSYS_UNCONNECTED__593, 
        SYNOPSYS_UNCONNECTED__594, SYNOPSYS_UNCONNECTED__595, 
        SYNOPSYS_UNCONNECTED__596, SYNOPSYS_UNCONNECTED__597, 
        SYNOPSYS_UNCONNECTED__598, SYNOPSYS_UNCONNECTED__599, 
        SYNOPSYS_UNCONNECTED__600, SYNOPSYS_UNCONNECTED__601, 
        SYNOPSYS_UNCONNECTED__602, SYNOPSYS_UNCONNECTED__603, 
        SYNOPSYS_UNCONNECTED__604, SYNOPSYS_UNCONNECTED__605, 
        SYNOPSYS_UNCONNECTED__606, SYNOPSYS_UNCONNECTED__607, 
        SYNOPSYS_UNCONNECTED__608, SYNOPSYS_UNCONNECTED__609, 
        SYNOPSYS_UNCONNECTED__610, SYNOPSYS_UNCONNECTED__611, 
        SYNOPSYS_UNCONNECTED__612, SYNOPSYS_UNCONNECTED__613, 
        SYNOPSYS_UNCONNECTED__614, SYNOPSYS_UNCONNECTED__615, 
        SYNOPSYS_UNCONNECTED__616, SYNOPSYS_UNCONNECTED__617, 
        SYNOPSYS_UNCONNECTED__618, SYNOPSYS_UNCONNECTED__619, 
        SYNOPSYS_UNCONNECTED__620, SYNOPSYS_UNCONNECTED__621, 
        SYNOPSYS_UNCONNECTED__622, SYNOPSYS_UNCONNECTED__623, 
        SYNOPSYS_UNCONNECTED__624, SYNOPSYS_UNCONNECTED__625, 
        SYNOPSYS_UNCONNECTED__626, SYNOPSYS_UNCONNECTED__627, 
        SYNOPSYS_UNCONNECTED__628, SYNOPSYS_UNCONNECTED__629, 
        SYNOPSYS_UNCONNECTED__630, SYNOPSYS_UNCONNECTED__631, 
        SYNOPSYS_UNCONNECTED__632, SYNOPSYS_UNCONNECTED__633, 
        SYNOPSYS_UNCONNECTED__634, SYNOPSYS_UNCONNECTED__635, 
        SYNOPSYS_UNCONNECTED__636, SYNOPSYS_UNCONNECTED__637, 
        SYNOPSYS_UNCONNECTED__638, SYNOPSYS_UNCONNECTED__639, 
        SYNOPSYS_UNCONNECTED__640, SYNOPSYS_UNCONNECTED__641, 
        SYNOPSYS_UNCONNECTED__642, SYNOPSYS_UNCONNECTED__643, 
        SYNOPSYS_UNCONNECTED__644, SYNOPSYS_UNCONNECTED__645, 
        SYNOPSYS_UNCONNECTED__646, SYNOPSYS_UNCONNECTED__647, 
        SYNOPSYS_UNCONNECTED__648, SYNOPSYS_UNCONNECTED__649, 
        SYNOPSYS_UNCONNECTED__650, SYNOPSYS_UNCONNECTED__651, 
        SYNOPSYS_UNCONNECTED__652, SYNOPSYS_UNCONNECTED__653, 
        SYNOPSYS_UNCONNECTED__654, SYNOPSYS_UNCONNECTED__655, 
        SYNOPSYS_UNCONNECTED__656, SYNOPSYS_UNCONNECTED__657, 
        SYNOPSYS_UNCONNECTED__658, SYNOPSYS_UNCONNECTED__659, 
        SYNOPSYS_UNCONNECTED__660, SYNOPSYS_UNCONNECTED__661, 
        SYNOPSYS_UNCONNECTED__662, SYNOPSYS_UNCONNECTED__663, 
        SYNOPSYS_UNCONNECTED__664, SYNOPSYS_UNCONNECTED__665, 
        SYNOPSYS_UNCONNECTED__666, SYNOPSYS_UNCONNECTED__667, 
        SYNOPSYS_UNCONNECTED__668, SYNOPSYS_UNCONNECTED__669, 
        SYNOPSYS_UNCONNECTED__670, SYNOPSYS_UNCONNECTED__671, 
        SYNOPSYS_UNCONNECTED__672, SYNOPSYS_UNCONNECTED__673, 
        SYNOPSYS_UNCONNECTED__674, SYNOPSYS_UNCONNECTED__675, 
        SYNOPSYS_UNCONNECTED__676, SYNOPSYS_UNCONNECTED__677, 
        SYNOPSYS_UNCONNECTED__678, SYNOPSYS_UNCONNECTED__679, 
        SYNOPSYS_UNCONNECTED__680, SYNOPSYS_UNCONNECTED__681, 
        SYNOPSYS_UNCONNECTED__682, SYNOPSYS_UNCONNECTED__683, 
        SYNOPSYS_UNCONNECTED__684, SYNOPSYS_UNCONNECTED__685, 
        SYNOPSYS_UNCONNECTED__686, SYNOPSYS_UNCONNECTED__687, 
        SYNOPSYS_UNCONNECTED__688, SYNOPSYS_UNCONNECTED__689, 
        SYNOPSYS_UNCONNECTED__690, SYNOPSYS_UNCONNECTED__691, 
        SYNOPSYS_UNCONNECTED__692, SYNOPSYS_UNCONNECTED__693, 
        SYNOPSYS_UNCONNECTED__694, SYNOPSYS_UNCONNECTED__695, 
        SYNOPSYS_UNCONNECTED__696, SYNOPSYS_UNCONNECTED__697, 
        SYNOPSYS_UNCONNECTED__698, SYNOPSYS_UNCONNECTED__699, 
        SYNOPSYS_UNCONNECTED__700, SYNOPSYS_UNCONNECTED__701, 
        SYNOPSYS_UNCONNECTED__702, SYNOPSYS_UNCONNECTED__703, 
        SYNOPSYS_UNCONNECTED__704, SYNOPSYS_UNCONNECTED__705, 
        SYNOPSYS_UNCONNECTED__706, SYNOPSYS_UNCONNECTED__707, 
        SYNOPSYS_UNCONNECTED__708, SYNOPSYS_UNCONNECTED__709, 
        SYNOPSYS_UNCONNECTED__710, SYNOPSYS_UNCONNECTED__711, 
        SYNOPSYS_UNCONNECTED__712, SYNOPSYS_UNCONNECTED__713, 
        SYNOPSYS_UNCONNECTED__714, SYNOPSYS_UNCONNECTED__715, 
        SYNOPSYS_UNCONNECTED__716, SYNOPSYS_UNCONNECTED__717, 
        SYNOPSYS_UNCONNECTED__718, SYNOPSYS_UNCONNECTED__719, 
        SYNOPSYS_UNCONNECTED__720, SYNOPSYS_UNCONNECTED__721, 
        SYNOPSYS_UNCONNECTED__722, SYNOPSYS_UNCONNECTED__723, 
        SYNOPSYS_UNCONNECTED__724, SYNOPSYS_UNCONNECTED__725, 
        SYNOPSYS_UNCONNECTED__726, SYNOPSYS_UNCONNECTED__727, 
        SYNOPSYS_UNCONNECTED__728, SYNOPSYS_UNCONNECTED__729, 
        SYNOPSYS_UNCONNECTED__730, SYNOPSYS_UNCONNECTED__731, 
        SYNOPSYS_UNCONNECTED__732, SYNOPSYS_UNCONNECTED__733, 
        SYNOPSYS_UNCONNECTED__734, SYNOPSYS_UNCONNECTED__735, 
        SYNOPSYS_UNCONNECTED__736, SYNOPSYS_UNCONNECTED__737, 
        SYNOPSYS_UNCONNECTED__738, SYNOPSYS_UNCONNECTED__739, 
        SYNOPSYS_UNCONNECTED__740, SYNOPSYS_UNCONNECTED__741, 
        SYNOPSYS_UNCONNECTED__742, SYNOPSYS_UNCONNECTED__743, 
        SYNOPSYS_UNCONNECTED__744, SYNOPSYS_UNCONNECTED__745, 
        SYNOPSYS_UNCONNECTED__746, SYNOPSYS_UNCONNECTED__747, 
        SYNOPSYS_UNCONNECTED__748, SYNOPSYS_UNCONNECTED__749, 
        SYNOPSYS_UNCONNECTED__750, SYNOPSYS_UNCONNECTED__751, 
        SYNOPSYS_UNCONNECTED__752, SYNOPSYS_UNCONNECTED__753, 
        SYNOPSYS_UNCONNECTED__754, SYNOPSYS_UNCONNECTED__755, 
        SYNOPSYS_UNCONNECTED__756, SYNOPSYS_UNCONNECTED__757, 
        SYNOPSYS_UNCONNECTED__758, SYNOPSYS_UNCONNECTED__759, 
        SYNOPSYS_UNCONNECTED__760, SYNOPSYS_UNCONNECTED__761, 
        SYNOPSYS_UNCONNECTED__762, SYNOPSYS_UNCONNECTED__763, 
        SYNOPSYS_UNCONNECTED__764, SYNOPSYS_UNCONNECTED__765, 
        SYNOPSYS_UNCONNECTED__766, SYNOPSYS_UNCONNECTED__767, 
        SYNOPSYS_UNCONNECTED__768, SYNOPSYS_UNCONNECTED__769, 
        SYNOPSYS_UNCONNECTED__770, SYNOPSYS_UNCONNECTED__771, 
        SYNOPSYS_UNCONNECTED__772, SYNOPSYS_UNCONNECTED__773, 
        SYNOPSYS_UNCONNECTED__774, SYNOPSYS_UNCONNECTED__775, 
        SYNOPSYS_UNCONNECTED__776, SYNOPSYS_UNCONNECTED__777, 
        SYNOPSYS_UNCONNECTED__778, SYNOPSYS_UNCONNECTED__779, 
        SYNOPSYS_UNCONNECTED__780, SYNOPSYS_UNCONNECTED__781, 
        SYNOPSYS_UNCONNECTED__782, SYNOPSYS_UNCONNECTED__783, 
        SYNOPSYS_UNCONNECTED__784, SYNOPSYS_UNCONNECTED__785, 
        SYNOPSYS_UNCONNECTED__786, SYNOPSYS_UNCONNECTED__787, 
        SYNOPSYS_UNCONNECTED__788, SYNOPSYS_UNCONNECTED__789, 
        SYNOPSYS_UNCONNECTED__790, SYNOPSYS_UNCONNECTED__791, 
        SYNOPSYS_UNCONNECTED__792, SYNOPSYS_UNCONNECTED__793, 
        SYNOPSYS_UNCONNECTED__794, SYNOPSYS_UNCONNECTED__795, 
        SYNOPSYS_UNCONNECTED__796, SYNOPSYS_UNCONNECTED__797, 
        SYNOPSYS_UNCONNECTED__798, SYNOPSYS_UNCONNECTED__799, 
        SYNOPSYS_UNCONNECTED__800, SYNOPSYS_UNCONNECTED__801, 
        SYNOPSYS_UNCONNECTED__802, SYNOPSYS_UNCONNECTED__803, 
        SYNOPSYS_UNCONNECTED__804, SYNOPSYS_UNCONNECTED__805, 
        SYNOPSYS_UNCONNECTED__806, SYNOPSYS_UNCONNECTED__807, 
        SYNOPSYS_UNCONNECTED__808, SYNOPSYS_UNCONNECTED__809, 
        SYNOPSYS_UNCONNECTED__810, SYNOPSYS_UNCONNECTED__811, 
        SYNOPSYS_UNCONNECTED__812, SYNOPSYS_UNCONNECTED__813, 
        SYNOPSYS_UNCONNECTED__814, SYNOPSYS_UNCONNECTED__815, 
        SYNOPSYS_UNCONNECTED__816, SYNOPSYS_UNCONNECTED__817, 
        SYNOPSYS_UNCONNECTED__818, SYNOPSYS_UNCONNECTED__819, 
        SYNOPSYS_UNCONNECTED__820, SYNOPSYS_UNCONNECTED__821, 
        SYNOPSYS_UNCONNECTED__822, SYNOPSYS_UNCONNECTED__823, 
        SYNOPSYS_UNCONNECTED__824, SYNOPSYS_UNCONNECTED__825, 
        SYNOPSYS_UNCONNECTED__826, SYNOPSYS_UNCONNECTED__827, 
        SYNOPSYS_UNCONNECTED__828, SYNOPSYS_UNCONNECTED__829, 
        SYNOPSYS_UNCONNECTED__830, SYNOPSYS_UNCONNECTED__831, 
        SYNOPSYS_UNCONNECTED__832, SYNOPSYS_UNCONNECTED__833, 
        SYNOPSYS_UNCONNECTED__834, SYNOPSYS_UNCONNECTED__835, 
        SYNOPSYS_UNCONNECTED__836, SYNOPSYS_UNCONNECTED__837, 
        SYNOPSYS_UNCONNECTED__838, SYNOPSYS_UNCONNECTED__839, 
        SYNOPSYS_UNCONNECTED__840, SYNOPSYS_UNCONNECTED__841, 
        SYNOPSYS_UNCONNECTED__842, SYNOPSYS_UNCONNECTED__843, 
        SYNOPSYS_UNCONNECTED__844, SYNOPSYS_UNCONNECTED__845, 
        SYNOPSYS_UNCONNECTED__846, SYNOPSYS_UNCONNECTED__847, 
        SYNOPSYS_UNCONNECTED__848, SYNOPSYS_UNCONNECTED__849, 
        SYNOPSYS_UNCONNECTED__850, SYNOPSYS_UNCONNECTED__851, 
        SYNOPSYS_UNCONNECTED__852, SYNOPSYS_UNCONNECTED__853, 
        SYNOPSYS_UNCONNECTED__854, SYNOPSYS_UNCONNECTED__855, 
        SYNOPSYS_UNCONNECTED__856, SYNOPSYS_UNCONNECTED__857, 
        SYNOPSYS_UNCONNECTED__858, SYNOPSYS_UNCONNECTED__859, 
        SYNOPSYS_UNCONNECTED__860, SYNOPSYS_UNCONNECTED__861, 
        SYNOPSYS_UNCONNECTED__862, SYNOPSYS_UNCONNECTED__863, 
        SYNOPSYS_UNCONNECTED__864, SYNOPSYS_UNCONNECTED__865, 
        SYNOPSYS_UNCONNECTED__866, SYNOPSYS_UNCONNECTED__867, 
        SYNOPSYS_UNCONNECTED__868, SYNOPSYS_UNCONNECTED__869, 
        SYNOPSYS_UNCONNECTED__870, SYNOPSYS_UNCONNECTED__871, 
        SYNOPSYS_UNCONNECTED__872, SYNOPSYS_UNCONNECTED__873, 
        SYNOPSYS_UNCONNECTED__874, SYNOPSYS_UNCONNECTED__875, 
        SYNOPSYS_UNCONNECTED__876, SYNOPSYS_UNCONNECTED__877, 
        SYNOPSYS_UNCONNECTED__878, SYNOPSYS_UNCONNECTED__879, 
        SYNOPSYS_UNCONNECTED__880, SYNOPSYS_UNCONNECTED__881, 
        SYNOPSYS_UNCONNECTED__882, SYNOPSYS_UNCONNECTED__883, 
        SYNOPSYS_UNCONNECTED__884, SYNOPSYS_UNCONNECTED__885, 
        SYNOPSYS_UNCONNECTED__886, SYNOPSYS_UNCONNECTED__887, 
        SYNOPSYS_UNCONNECTED__888, SYNOPSYS_UNCONNECTED__889, 
        SYNOPSYS_UNCONNECTED__890, SYNOPSYS_UNCONNECTED__891, 
        SYNOPSYS_UNCONNECTED__892, SYNOPSYS_UNCONNECTED__893, 
        SYNOPSYS_UNCONNECTED__894, SYNOPSYS_UNCONNECTED__895, 
        SYNOPSYS_UNCONNECTED__896, SYNOPSYS_UNCONNECTED__897, 
        SYNOPSYS_UNCONNECTED__898, SYNOPSYS_UNCONNECTED__899, 
        SYNOPSYS_UNCONNECTED__900, SYNOPSYS_UNCONNECTED__901, 
        SYNOPSYS_UNCONNECTED__902, SYNOPSYS_UNCONNECTED__903, 
        SYNOPSYS_UNCONNECTED__904, SYNOPSYS_UNCONNECTED__905, 
        SYNOPSYS_UNCONNECTED__906, SYNOPSYS_UNCONNECTED__907, 
        SYNOPSYS_UNCONNECTED__908, SYNOPSYS_UNCONNECTED__909, 
        SYNOPSYS_UNCONNECTED__910, SYNOPSYS_UNCONNECTED__911, 
        SYNOPSYS_UNCONNECTED__912, SYNOPSYS_UNCONNECTED__913, 
        SYNOPSYS_UNCONNECTED__914, SYNOPSYS_UNCONNECTED__915, 
        SYNOPSYS_UNCONNECTED__916, SYNOPSYS_UNCONNECTED__917, 
        SYNOPSYS_UNCONNECTED__918, SYNOPSYS_UNCONNECTED__919, 
        SYNOPSYS_UNCONNECTED__920, SYNOPSYS_UNCONNECTED__921, 
        SYNOPSYS_UNCONNECTED__922, SYNOPSYS_UNCONNECTED__923, 
        SYNOPSYS_UNCONNECTED__924, SYNOPSYS_UNCONNECTED__925, 
        SYNOPSYS_UNCONNECTED__926, SYNOPSYS_UNCONNECTED__927, 
        SYNOPSYS_UNCONNECTED__928, SYNOPSYS_UNCONNECTED__929, 
        SYNOPSYS_UNCONNECTED__930, SYNOPSYS_UNCONNECTED__931, 
        SYNOPSYS_UNCONNECTED__932, SYNOPSYS_UNCONNECTED__933, 
        SYNOPSYS_UNCONNECTED__934, SYNOPSYS_UNCONNECTED__935, 
        SYNOPSYS_UNCONNECTED__936, SYNOPSYS_UNCONNECTED__937, 
        SYNOPSYS_UNCONNECTED__938, SYNOPSYS_UNCONNECTED__939, 
        SYNOPSYS_UNCONNECTED__940, SYNOPSYS_UNCONNECTED__941, 
        SYNOPSYS_UNCONNECTED__942, SYNOPSYS_UNCONNECTED__943, 
        SYNOPSYS_UNCONNECTED__944, SYNOPSYS_UNCONNECTED__945, 
        SYNOPSYS_UNCONNECTED__946, SYNOPSYS_UNCONNECTED__947, 
        SYNOPSYS_UNCONNECTED__948, SYNOPSYS_UNCONNECTED__949, 
        SYNOPSYS_UNCONNECTED__950, SYNOPSYS_UNCONNECTED__951, 
        SYNOPSYS_UNCONNECTED__952, SYNOPSYS_UNCONNECTED__953, 
        SYNOPSYS_UNCONNECTED__954, SYNOPSYS_UNCONNECTED__955, 
        SYNOPSYS_UNCONNECTED__956, SYNOPSYS_UNCONNECTED__957, 
        SYNOPSYS_UNCONNECTED__958, SYNOPSYS_UNCONNECTED__959, 
        SYNOPSYS_UNCONNECTED__960, SYNOPSYS_UNCONNECTED__961, 
        SYNOPSYS_UNCONNECTED__962, SYNOPSYS_UNCONNECTED__963, 
        SYNOPSYS_UNCONNECTED__964, SYNOPSYS_UNCONNECTED__965, 
        SYNOPSYS_UNCONNECTED__966, SYNOPSYS_UNCONNECTED__967, 
        SYNOPSYS_UNCONNECTED__968, SYNOPSYS_UNCONNECTED__969, 
        SYNOPSYS_UNCONNECTED__970, SYNOPSYS_UNCONNECTED__971, 
        SYNOPSYS_UNCONNECTED__972, SYNOPSYS_UNCONNECTED__973, 
        SYNOPSYS_UNCONNECTED__974, SYNOPSYS_UNCONNECTED__975, 
        SYNOPSYS_UNCONNECTED__976, SYNOPSYS_UNCONNECTED__977, 
        SYNOPSYS_UNCONNECTED__978, SYNOPSYS_UNCONNECTED__979, 
        SYNOPSYS_UNCONNECTED__980, SYNOPSYS_UNCONNECTED__981, 
        SYNOPSYS_UNCONNECTED__982, SYNOPSYS_UNCONNECTED__983, 
        SYNOPSYS_UNCONNECTED__984, SYNOPSYS_UNCONNECTED__985, 
        SYNOPSYS_UNCONNECTED__986, SYNOPSYS_UNCONNECTED__987, 
        SYNOPSYS_UNCONNECTED__988, SYNOPSYS_UNCONNECTED__989, 
        SYNOPSYS_UNCONNECTED__990, SYNOPSYS_UNCONNECTED__991, 
        SYNOPSYS_UNCONNECTED__992, SYNOPSYS_UNCONNECTED__993, 
        SYNOPSYS_UNCONNECTED__994, SYNOPSYS_UNCONNECTED__995, 
        SYNOPSYS_UNCONNECTED__996, SYNOPSYS_UNCONNECTED__997, 
        SYNOPSYS_UNCONNECTED__998, SYNOPSYS_UNCONNECTED__999, 
        SYNOPSYS_UNCONNECTED__1000, SYNOPSYS_UNCONNECTED__1001, 
        SYNOPSYS_UNCONNECTED__1002, SYNOPSYS_UNCONNECTED__1003, 
        SYNOPSYS_UNCONNECTED__1004, SYNOPSYS_UNCONNECTED__1005, 
        SYNOPSYS_UNCONNECTED__1006, SYNOPSYS_UNCONNECTED__1007, 
        SYNOPSYS_UNCONNECTED__1008, SYNOPSYS_UNCONNECTED__1009, 
        SYNOPSYS_UNCONNECTED__1010, SYNOPSYS_UNCONNECTED__1011, 
        SYNOPSYS_UNCONNECTED__1012, SYNOPSYS_UNCONNECTED__1013, 
        SYNOPSYS_UNCONNECTED__1014, SYNOPSYS_UNCONNECTED__1015, 
        SYNOPSYS_UNCONNECTED__1016, SYNOPSYS_UNCONNECTED__1017, 
        SYNOPSYS_UNCONNECTED__1018, SYNOPSYS_UNCONNECTED__1019, 
        SYNOPSYS_UNCONNECTED__1020, SYNOPSYS_UNCONNECTED__1021, 
        SYNOPSYS_UNCONNECTED__1022, SYNOPSYS_UNCONNECTED__1023, 
        SYNOPSYS_UNCONNECTED__1024, SYNOPSYS_UNCONNECTED__1025, 
        SYNOPSYS_UNCONNECTED__1026, SYNOPSYS_UNCONNECTED__1027, 
        SYNOPSYS_UNCONNECTED__1028, SYNOPSYS_UNCONNECTED__1029, 
        SYNOPSYS_UNCONNECTED__1030, SYNOPSYS_UNCONNECTED__1031, 
        SYNOPSYS_UNCONNECTED__1032, SYNOPSYS_UNCONNECTED__1033, 
        SYNOPSYS_UNCONNECTED__1034, SYNOPSYS_UNCONNECTED__1035, 
        SYNOPSYS_UNCONNECTED__1036, SYNOPSYS_UNCONNECTED__1037, 
        SYNOPSYS_UNCONNECTED__1038, SYNOPSYS_UNCONNECTED__1039, 
        SYNOPSYS_UNCONNECTED__1040, SYNOPSYS_UNCONNECTED__1041, 
        SYNOPSYS_UNCONNECTED__1042, SYNOPSYS_UNCONNECTED__1043, 
        SYNOPSYS_UNCONNECTED__1044, SYNOPSYS_UNCONNECTED__1045, 
        SYNOPSYS_UNCONNECTED__1046, SYNOPSYS_UNCONNECTED__1047, 
        SYNOPSYS_UNCONNECTED__1048, SYNOPSYS_UNCONNECTED__1049, 
        SYNOPSYS_UNCONNECTED__1050, SYNOPSYS_UNCONNECTED__1051, 
        SYNOPSYS_UNCONNECTED__1052, SYNOPSYS_UNCONNECTED__1053, 
        SYNOPSYS_UNCONNECTED__1054, SYNOPSYS_UNCONNECTED__1055, 
        SYNOPSYS_UNCONNECTED__1056, SYNOPSYS_UNCONNECTED__1057, 
        SYNOPSYS_UNCONNECTED__1058, SYNOPSYS_UNCONNECTED__1059, 
        SYNOPSYS_UNCONNECTED__1060, SYNOPSYS_UNCONNECTED__1061, 
        SYNOPSYS_UNCONNECTED__1062, SYNOPSYS_UNCONNECTED__1063, 
        SYNOPSYS_UNCONNECTED__1064, SYNOPSYS_UNCONNECTED__1065, 
        SYNOPSYS_UNCONNECTED__1066, SYNOPSYS_UNCONNECTED__1067, 
        SYNOPSYS_UNCONNECTED__1068, SYNOPSYS_UNCONNECTED__1069, 
        SYNOPSYS_UNCONNECTED__1070, SYNOPSYS_UNCONNECTED__1071, 
        SYNOPSYS_UNCONNECTED__1072, SYNOPSYS_UNCONNECTED__1073, 
        SYNOPSYS_UNCONNECTED__1074, SYNOPSYS_UNCONNECTED__1075, 
        SYNOPSYS_UNCONNECTED__1076, SYNOPSYS_UNCONNECTED__1077, 
        SYNOPSYS_UNCONNECTED__1078, SYNOPSYS_UNCONNECTED__1079, 
        SYNOPSYS_UNCONNECTED__1080, SYNOPSYS_UNCONNECTED__1081, 
        SYNOPSYS_UNCONNECTED__1082, SYNOPSYS_UNCONNECTED__1083, 
        SYNOPSYS_UNCONNECTED__1084, SYNOPSYS_UNCONNECTED__1085, 
        SYNOPSYS_UNCONNECTED__1086, SYNOPSYS_UNCONNECTED__1087, 
        SYNOPSYS_UNCONNECTED__1088, SYNOPSYS_UNCONNECTED__1089, 
        SYNOPSYS_UNCONNECTED__1090, SYNOPSYS_UNCONNECTED__1091, 
        SYNOPSYS_UNCONNECTED__1092, SYNOPSYS_UNCONNECTED__1093, 
        SYNOPSYS_UNCONNECTED__1094, SYNOPSYS_UNCONNECTED__1095, 
        SYNOPSYS_UNCONNECTED__1096, SYNOPSYS_UNCONNECTED__1097, 
        SYNOPSYS_UNCONNECTED__1098, SYNOPSYS_UNCONNECTED__1099, 
        SYNOPSYS_UNCONNECTED__1100, SYNOPSYS_UNCONNECTED__1101, 
        SYNOPSYS_UNCONNECTED__1102, SYNOPSYS_UNCONNECTED__1103, 
        SYNOPSYS_UNCONNECTED__1104, SYNOPSYS_UNCONNECTED__1105, 
        SYNOPSYS_UNCONNECTED__1106, SYNOPSYS_UNCONNECTED__1107, 
        SYNOPSYS_UNCONNECTED__1108, SYNOPSYS_UNCONNECTED__1109, 
        SYNOPSYS_UNCONNECTED__1110, SYNOPSYS_UNCONNECTED__1111, 
        SYNOPSYS_UNCONNECTED__1112, SYNOPSYS_UNCONNECTED__1113, 
        SYNOPSYS_UNCONNECTED__1114, SYNOPSYS_UNCONNECTED__1115, 
        SYNOPSYS_UNCONNECTED__1116, SYNOPSYS_UNCONNECTED__1117, 
        SYNOPSYS_UNCONNECTED__1118, SYNOPSYS_UNCONNECTED__1119, 
        SYNOPSYS_UNCONNECTED__1120, SYNOPSYS_UNCONNECTED__1121, 
        SYNOPSYS_UNCONNECTED__1122, SYNOPSYS_UNCONNECTED__1123, 
        SYNOPSYS_UNCONNECTED__1124, SYNOPSYS_UNCONNECTED__1125, 
        SYNOPSYS_UNCONNECTED__1126, SYNOPSYS_UNCONNECTED__1127, 
        SYNOPSYS_UNCONNECTED__1128, SYNOPSYS_UNCONNECTED__1129, 
        SYNOPSYS_UNCONNECTED__1130, SYNOPSYS_UNCONNECTED__1131, 
        SYNOPSYS_UNCONNECTED__1132, SYNOPSYS_UNCONNECTED__1133, 
        SYNOPSYS_UNCONNECTED__1134, SYNOPSYS_UNCONNECTED__1135, 
        SYNOPSYS_UNCONNECTED__1136, SYNOPSYS_UNCONNECTED__1137, 
        SYNOPSYS_UNCONNECTED__1138, SYNOPSYS_UNCONNECTED__1139, 
        SYNOPSYS_UNCONNECTED__1140, SYNOPSYS_UNCONNECTED__1141, 
        SYNOPSYS_UNCONNECTED__1142, SYNOPSYS_UNCONNECTED__1143, 
        SYNOPSYS_UNCONNECTED__1144, SYNOPSYS_UNCONNECTED__1145, 
        SYNOPSYS_UNCONNECTED__1146, SYNOPSYS_UNCONNECTED__1147, 
        SYNOPSYS_UNCONNECTED__1148, SYNOPSYS_UNCONNECTED__1149, 
        SYNOPSYS_UNCONNECTED__1150, SYNOPSYS_UNCONNECTED__1151, 
        SYNOPSYS_UNCONNECTED__1152, SYNOPSYS_UNCONNECTED__1153, 
        SYNOPSYS_UNCONNECTED__1154, SYNOPSYS_UNCONNECTED__1155, 
        SYNOPSYS_UNCONNECTED__1156, SYNOPSYS_UNCONNECTED__1157, 
        SYNOPSYS_UNCONNECTED__1158, SYNOPSYS_UNCONNECTED__1159, 
        SYNOPSYS_UNCONNECTED__1160, SYNOPSYS_UNCONNECTED__1161, 
        SYNOPSYS_UNCONNECTED__1162, SYNOPSYS_UNCONNECTED__1163, 
        SYNOPSYS_UNCONNECTED__1164, SYNOPSYS_UNCONNECTED__1165, 
        SYNOPSYS_UNCONNECTED__1166, SYNOPSYS_UNCONNECTED__1167, 
        SYNOPSYS_UNCONNECTED__1168, SYNOPSYS_UNCONNECTED__1169, 
        SYNOPSYS_UNCONNECTED__1170, SYNOPSYS_UNCONNECTED__1171, 
        SYNOPSYS_UNCONNECTED__1172, SYNOPSYS_UNCONNECTED__1173, 
        SYNOPSYS_UNCONNECTED__1174, SYNOPSYS_UNCONNECTED__1175, 
        SYNOPSYS_UNCONNECTED__1176, SYNOPSYS_UNCONNECTED__1177, 
        SYNOPSYS_UNCONNECTED__1178, SYNOPSYS_UNCONNECTED__1179, 
        SYNOPSYS_UNCONNECTED__1180, SYNOPSYS_UNCONNECTED__1181, 
        SYNOPSYS_UNCONNECTED__1182, SYNOPSYS_UNCONNECTED__1183, 
        SYNOPSYS_UNCONNECTED__1184, SYNOPSYS_UNCONNECTED__1185, 
        SYNOPSYS_UNCONNECTED__1186, SYNOPSYS_UNCONNECTED__1187, 
        SYNOPSYS_UNCONNECTED__1188, SYNOPSYS_UNCONNECTED__1189, 
        SYNOPSYS_UNCONNECTED__1190, SYNOPSYS_UNCONNECTED__1191, 
        SYNOPSYS_UNCONNECTED__1192, SYNOPSYS_UNCONNECTED__1193, 
        SYNOPSYS_UNCONNECTED__1194, SYNOPSYS_UNCONNECTED__1195, 
        SYNOPSYS_UNCONNECTED__1196, SYNOPSYS_UNCONNECTED__1197, 
        SYNOPSYS_UNCONNECTED__1198, SYNOPSYS_UNCONNECTED__1199, 
        SYNOPSYS_UNCONNECTED__1200, SYNOPSYS_UNCONNECTED__1201, 
        SYNOPSYS_UNCONNECTED__1202, SYNOPSYS_UNCONNECTED__1203, 
        SYNOPSYS_UNCONNECTED__1204, SYNOPSYS_UNCONNECTED__1205, 
        SYNOPSYS_UNCONNECTED__1206, SYNOPSYS_UNCONNECTED__1207, 
        SYNOPSYS_UNCONNECTED__1208, SYNOPSYS_UNCONNECTED__1209, 
        SYNOPSYS_UNCONNECTED__1210, SYNOPSYS_UNCONNECTED__1211, 
        SYNOPSYS_UNCONNECTED__1212, SYNOPSYS_UNCONNECTED__1213, 
        SYNOPSYS_UNCONNECTED__1214, SYNOPSYS_UNCONNECTED__1215, 
        SYNOPSYS_UNCONNECTED__1216, SYNOPSYS_UNCONNECTED__1217, 
        SYNOPSYS_UNCONNECTED__1218, SYNOPSYS_UNCONNECTED__1219, 
        SYNOPSYS_UNCONNECTED__1220, SYNOPSYS_UNCONNECTED__1221, 
        SYNOPSYS_UNCONNECTED__1222, SYNOPSYS_UNCONNECTED__1223, 
        SYNOPSYS_UNCONNECTED__1224, SYNOPSYS_UNCONNECTED__1225, 
        SYNOPSYS_UNCONNECTED__1226, SYNOPSYS_UNCONNECTED__1227, 
        SYNOPSYS_UNCONNECTED__1228, SYNOPSYS_UNCONNECTED__1229, 
        SYNOPSYS_UNCONNECTED__1230, SYNOPSYS_UNCONNECTED__1231;

  ADDER_P4_N_BIT64_0 adder_1 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, \mux_out[1][31] , \mux_out[1][30] , \mux_out[1][29] , 
        \mux_out[1][28] , \mux_out[1][27] , \mux_out[1][26] , \mux_out[1][25] , 
        \mux_out[1][24] , \mux_out[1][23] , \mux_out[1][22] , \mux_out[1][21] , 
        \mux_out[1][20] , \mux_out[1][19] , \mux_out[1][18] , \mux_out[1][17] , 
        \mux_out[1][16] , \mux_out[1][15] , \mux_out[1][14] , \mux_out[1][13] , 
        \mux_out[1][12] , \mux_out[1][11] , \mux_out[1][10] , \mux_out[1][9] , 
        \mux_out[1][8] , \mux_out[1][7] , \mux_out[1][6] , \mux_out[1][5] , 
        \mux_out[1][4] , \mux_out[1][3] , \mux_out[1][2] , 1'b0, 1'b0}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \add_out_s1[0][31] , 
        \add_out_s1[0][30] , \add_out_s1[0][29] , \add_out_s1[0][28] , 
        \add_out_s1[0][27] , \add_out_s1[0][26] , \add_out_s1[0][25] , 
        \add_out_s1[0][24] , \add_out_s1[0][23] , \add_out_s1[0][22] , 
        \add_out_s1[0][21] , \add_out_s1[0][20] , \add_out_s1[0][19] , 
        \add_out_s1[0][18] , \add_out_s1[0][17] , \add_out_s1[0][16] , 
        \add_out_s1[0][15] , \add_out_s1[0][14] , \add_out_s1[0][13] , 
        \add_out_s1[0][12] , \add_out_s1[0][11] , \add_out_s1[0][10] , 
        \add_out_s1[0][9] , \add_out_s1[0][8] , \add_out_s1[0][7] , 
        \add_out_s1[0][6] , \add_out_s1[0][5] , \add_out_s1[0][4] , 
        \add_out_s1[0][3] , \add_out_s1[0][2] , \add_out_s1[0][1] , 
        \add_out_s1[0][0] }), .add_sub(1'b0), .SUM({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, SYNOPSYS_UNCONNECTED__22, 
        SYNOPSYS_UNCONNECTED__23, SYNOPSYS_UNCONNECTED__24, 
        SYNOPSYS_UNCONNECTED__25, SYNOPSYS_UNCONNECTED__26, 
        SYNOPSYS_UNCONNECTED__27, SYNOPSYS_UNCONNECTED__28, 
        SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, 
        SYNOPSYS_UNCONNECTED__31, \add_out_s1[1][31] , \add_out_s1[1][30] , 
        \add_out_s1[1][29] , \add_out_s1[1][28] , \add_out_s1[1][27] , 
        \add_out_s1[1][26] , \add_out_s1[1][25] , n16, \add_out_s1[1][23] , 
        \add_out_s1[1][22] , \add_out_s1[1][21] , \add_out_s1[1][20] , 
        \add_out_s1[1][19] , \add_out_s1[1][18] , \add_out_s1[1][17] , 
        \add_out_s1[1][16] , \add_out_s1[1][15] , \add_out_s1[1][14] , 
        \add_out_s1[1][13] , \add_out_s1[1][12] , \add_out_s1[1][11] , 
        \add_out_s1[1][10] , \add_out_s1[1][9] , \add_out_s1[1][8] , 
        \add_out_s1[1][7] , \add_out_s1[1][6] , \add_out_s1[1][5] , 
        \add_out_s1[1][4] , \add_out_s1[1][3] , \add_out_s1[1][2] , 
        \add_out_s1[1][1] , \add_out_s1[1][0] }) );
  ADDER_P4_N_BIT64_14 adder_2 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, \mux_out[2][31] , \mux_out[2][30] , \mux_out[2][29] , 
        \mux_out[2][28] , \mux_out[2][27] , \mux_out[2][26] , \mux_out[2][25] , 
        \mux_out[2][24] , \mux_out[2][23] , \mux_out[2][22] , \mux_out[2][21] , 
        \mux_out[2][20] , \mux_out[2][19] , \mux_out[2][18] , \mux_out[2][17] , 
        \mux_out[2][16] , \mux_out[2][15] , \mux_out[2][14] , \mux_out[2][13] , 
        \mux_out[2][12] , \mux_out[2][11] , \mux_out[2][10] , \mux_out[2][9] , 
        \mux_out[2][8] , \mux_out[2][7] , \mux_out[2][6] , \mux_out[2][5] , 
        \mux_out[2][4] , 1'b0, 1'b0, 1'b0, 1'b0}), .B({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, \add_out_s1[1][31] , \add_out_s1[1][30] , 
        \add_out_s1[1][29] , \add_out_s1[1][28] , \add_out_s1[1][27] , 
        \add_out_s1[1][26] , \add_out_s1[1][25] , n16, \add_out_s1[1][23] , 
        \add_out_s1[1][22] , \add_out_s1[1][21] , \add_out_s1[1][20] , 
        \add_out_s1[1][19] , \add_out_s1[1][18] , \add_out_s1[1][17] , 
        \add_out_s1[1][16] , \add_out_s1[1][15] , \add_out_s1[1][14] , 
        \add_out_s1[1][13] , \add_out_s1[1][12] , \add_out_s1[1][11] , 
        \add_out_s1[1][10] , \add_out_s1[1][9] , \add_out_s1[1][8] , 
        \add_out_s1[1][7] , \add_out_s1[1][6] , \add_out_s1[1][5] , 
        \add_out_s1[1][4] , \add_out_s1[1][3] , \add_out_s1[1][2] , 
        \add_out_s1[1][1] , \add_out_s1[1][0] }), .add_sub(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        \add_out_s1[2][31] , \add_out_s1[2][30] , \add_out_s1[2][29] , 
        \add_out_s1[2][28] , \add_out_s1[2][27] , \add_out_s1[2][26] , 
        \add_out_s1[2][25] , \add_out_s1[2][24] , \add_out_s1[2][23] , 
        \add_out_s1[2][22] , \add_out_s1[2][21] , \add_out_s1[2][20] , 
        \add_out_s1[2][19] , \add_out_s1[2][18] , \add_out_s1[2][17] , 
        \add_out_s1[2][16] , \add_out_s1[2][15] , \add_out_s1[2][14] , 
        \add_out_s1[2][13] , \add_out_s1[2][12] , \add_out_s1[2][11] , 
        \add_out_s1[2][10] , \add_out_s1[2][9] , \add_out_s1[2][8] , 
        \add_out_s1[2][7] , \add_out_s1[2][6] , \add_out_s1[2][5] , 
        \add_out_s1[2][4] , \add_out_s1[2][3] , \add_out_s1[2][2] , 
        \add_out_s1[2][1] , \add_out_s1[2][0] }) );
  ADDER_P4_N_BIT64_13 adder_3 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, \mux_out[3][31] , \mux_out[3][30] , \mux_out[3][29] , 
        \mux_out[3][28] , \mux_out[3][27] , \mux_out[3][26] , \mux_out[3][25] , 
        \mux_out[3][24] , \mux_out[3][23] , \mux_out[3][22] , \mux_out[3][21] , 
        \mux_out[3][20] , \mux_out[3][19] , \mux_out[3][18] , \mux_out[3][17] , 
        \mux_out[3][16] , \mux_out[3][15] , \mux_out[3][14] , \mux_out[3][13] , 
        \mux_out[3][12] , \mux_out[3][11] , \mux_out[3][10] , \mux_out[3][9] , 
        \mux_out[3][8] , \mux_out[3][7] , \mux_out[3][6] , 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        \add_out_s1[2][31] , \add_out_s1[2][30] , \add_out_s1[2][29] , 
        \add_out_s1[2][28] , \add_out_s1[2][27] , \add_out_s1[2][26] , 
        \add_out_s1[2][25] , \add_out_s1[2][24] , \add_out_s1[2][23] , 
        \add_out_s1[2][22] , \add_out_s1[2][21] , \add_out_s1[2][20] , 
        \add_out_s1[2][19] , \add_out_s1[2][18] , \add_out_s1[2][17] , 
        \add_out_s1[2][16] , \add_out_s1[2][15] , \add_out_s1[2][14] , 
        \add_out_s1[2][13] , \add_out_s1[2][12] , \add_out_s1[2][11] , 
        \add_out_s1[2][10] , \add_out_s1[2][9] , \add_out_s1[2][8] , 
        \add_out_s1[2][7] , \add_out_s1[2][6] , \add_out_s1[2][5] , 
        \add_out_s1[2][4] , \add_out_s1[2][3] , \add_out_s1[2][2] , 
        \add_out_s1[2][1] , \add_out_s1[2][0] }), .add_sub(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        \add_out_s1[3][31] , \add_out_s1[3][30] , \add_out_s1[3][29] , 
        \add_out_s1[3][28] , \add_out_s1[3][27] , \add_out_s1[3][26] , 
        \add_out_s1[3][25] , \add_out_s1[3][24] , \add_out_s1[3][23] , 
        \add_out_s1[3][22] , \add_out_s1[3][21] , \add_out_s1[3][20] , 
        \add_out_s1[3][19] , \add_out_s1[3][18] , \add_out_s1[3][17] , 
        \add_out_s1[3][16] , n15, \add_out_s1[3][14] , \add_out_s1[3][13] , 
        \add_out_s1[3][12] , \add_out_s1[3][11] , \add_out_s1[3][10] , 
        \add_out_s1[3][9] , \add_out_s1[3][8] , \add_out_s1[3][7] , 
        \add_out_s1[3][6] , \add_out_s1[3][5] , \add_out_s1[3][4] , 
        \add_out_s1[3][3] , \add_out_s1[3][2] , \add_out_s1[3][1] , 
        \add_out_s1[3][0] }) );
  ADDER_P4_N_BIT64_12 adder_4 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, \mux_out[4][31] , \mux_out[4][30] , \mux_out[4][29] , 
        \mux_out[4][28] , \mux_out[4][27] , \mux_out[4][26] , \mux_out[4][25] , 
        \mux_out[4][24] , \mux_out[4][23] , \mux_out[4][22] , \mux_out[4][21] , 
        \mux_out[4][20] , \mux_out[4][19] , \mux_out[4][18] , \mux_out[4][17] , 
        \mux_out[4][16] , \mux_out[4][15] , \mux_out[4][14] , \mux_out[4][13] , 
        \mux_out[4][12] , \mux_out[4][11] , \mux_out[4][10] , \mux_out[4][9] , 
        \mux_out[4][8] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B(
        {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        \add_out_s1[3][31] , \add_out_s1[3][30] , \add_out_s1[3][29] , 
        \add_out_s1[3][28] , \add_out_s1[3][27] , \add_out_s1[3][26] , 
        \add_out_s1[3][25] , \add_out_s1[3][24] , \add_out_s1[3][23] , 
        \add_out_s1[3][22] , \add_out_s1[3][21] , \add_out_s1[3][20] , 
        \add_out_s1[3][19] , \add_out_s1[3][18] , \add_out_s1[3][17] , 
        \add_out_s1[3][16] , n15, \add_out_s1[3][14] , \add_out_s1[3][13] , 
        \add_out_s1[3][12] , \add_out_s1[3][11] , \add_out_s1[3][10] , 
        \add_out_s1[3][9] , \add_out_s1[3][8] , \add_out_s1[3][7] , 
        \add_out_s1[3][6] , \add_out_s1[3][5] , \add_out_s1[3][4] , 
        \add_out_s1[3][3] , \add_out_s1[3][2] , \add_out_s1[3][1] , 
        \add_out_s1[3][0] }), .add_sub(1'b0), .SUM({SYNOPSYS_UNCONNECTED__96, 
        SYNOPSYS_UNCONNECTED__97, SYNOPSYS_UNCONNECTED__98, 
        SYNOPSYS_UNCONNECTED__99, SYNOPSYS_UNCONNECTED__100, 
        SYNOPSYS_UNCONNECTED__101, SYNOPSYS_UNCONNECTED__102, 
        SYNOPSYS_UNCONNECTED__103, SYNOPSYS_UNCONNECTED__104, 
        SYNOPSYS_UNCONNECTED__105, SYNOPSYS_UNCONNECTED__106, 
        SYNOPSYS_UNCONNECTED__107, SYNOPSYS_UNCONNECTED__108, 
        SYNOPSYS_UNCONNECTED__109, SYNOPSYS_UNCONNECTED__110, 
        SYNOPSYS_UNCONNECTED__111, SYNOPSYS_UNCONNECTED__112, 
        SYNOPSYS_UNCONNECTED__113, SYNOPSYS_UNCONNECTED__114, 
        SYNOPSYS_UNCONNECTED__115, SYNOPSYS_UNCONNECTED__116, 
        SYNOPSYS_UNCONNECTED__117, SYNOPSYS_UNCONNECTED__118, 
        SYNOPSYS_UNCONNECTED__119, SYNOPSYS_UNCONNECTED__120, 
        SYNOPSYS_UNCONNECTED__121, SYNOPSYS_UNCONNECTED__122, 
        SYNOPSYS_UNCONNECTED__123, SYNOPSYS_UNCONNECTED__124, 
        SYNOPSYS_UNCONNECTED__125, SYNOPSYS_UNCONNECTED__126, 
        SYNOPSYS_UNCONNECTED__127, \add_out_s1[4][31] , \add_out_s1[4][30] , 
        \add_out_s1[4][29] , \add_out_s1[4][28] , \add_out_s1[4][27] , 
        \add_out_s1[4][26] , \add_out_s1[4][25] , \add_out_s1[4][24] , 
        \add_out_s1[4][23] , \add_out_s1[4][22] , \add_out_s1[4][21] , 
        \add_out_s1[4][20] , \add_out_s1[4][19] , \add_out_s1[4][18] , 
        \add_out_s1[4][17] , \add_out_s1[4][16] , \add_out_s1[4][15] , 
        \add_out_s1[4][14] , \add_out_s1[4][13] , \add_out_s1[4][12] , 
        \add_out_s1[4][11] , \add_out_s1[4][10] , \add_out_s1[4][9] , 
        \add_out_s1[4][8] , \add_out_s1[4][7] , \add_out_s1[4][6] , 
        \add_out_s1[4][5] , \add_out_s1[4][4] , \add_out_s1[4][3] , 
        \add_out_s1[4][2] , \add_out_s1[4][1] , \add_out_s1[4][0] }) );
  ADDER_P4_N_BIT64_11 adder_5 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, \mux_out[5][31] , \mux_out[5][30] , \mux_out[5][29] , 
        \mux_out[5][28] , \mux_out[5][27] , \mux_out[5][26] , \mux_out[5][25] , 
        \mux_out[5][24] , \mux_out[5][23] , \mux_out[5][22] , \mux_out[5][21] , 
        n22, \mux_out[5][19] , \mux_out[5][18] , \mux_out[5][17] , 
        \mux_out[5][16] , \mux_out[5][15] , \mux_out[5][14] , \mux_out[5][13] , 
        \mux_out[5][12] , \mux_out[5][11] , \mux_out[5][10] , 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, \add_out_s2[4][31] , \add_out_s2[4][30] , 
        \add_out_s2[4][29] , \add_out_s2[4][28] , \add_out_s2[4][27] , 
        \add_out_s2[4][26] , \add_out_s2[4][25] , \add_out_s2[4][24] , 
        \add_out_s2[4][23] , \add_out_s2[4][22] , \add_out_s2[4][21] , 
        \add_out_s2[4][20] , \add_out_s2[4][19] , \add_out_s2[4][18] , 
        \add_out_s2[4][17] , \add_out_s2[4][16] , \add_out_s2[4][15] , 
        \add_out_s2[4][14] , \add_out_s2[4][13] , \add_out_s2[4][12] , 
        \add_out_s2[4][11] , \add_out_s2[4][10] , \add_out_s2[4][9] , 
        \add_out_s2[4][8] , \add_out_s2[4][7] , \add_out_s2[4][6] , 
        \add_out_s2[4][5] , \add_out_s2[4][4] , \add_out_s2[4][3] , 
        \add_out_s2[4][2] , \add_out_s2[4][1] , \add_out_s2[4][0] }), 
        .add_sub(1'b0), .SUM({SYNOPSYS_UNCONNECTED__128, 
        SYNOPSYS_UNCONNECTED__129, SYNOPSYS_UNCONNECTED__130, 
        SYNOPSYS_UNCONNECTED__131, SYNOPSYS_UNCONNECTED__132, 
        SYNOPSYS_UNCONNECTED__133, SYNOPSYS_UNCONNECTED__134, 
        SYNOPSYS_UNCONNECTED__135, SYNOPSYS_UNCONNECTED__136, 
        SYNOPSYS_UNCONNECTED__137, SYNOPSYS_UNCONNECTED__138, 
        SYNOPSYS_UNCONNECTED__139, SYNOPSYS_UNCONNECTED__140, 
        SYNOPSYS_UNCONNECTED__141, SYNOPSYS_UNCONNECTED__142, 
        SYNOPSYS_UNCONNECTED__143, SYNOPSYS_UNCONNECTED__144, 
        SYNOPSYS_UNCONNECTED__145, SYNOPSYS_UNCONNECTED__146, 
        SYNOPSYS_UNCONNECTED__147, SYNOPSYS_UNCONNECTED__148, 
        SYNOPSYS_UNCONNECTED__149, SYNOPSYS_UNCONNECTED__150, 
        SYNOPSYS_UNCONNECTED__151, SYNOPSYS_UNCONNECTED__152, 
        SYNOPSYS_UNCONNECTED__153, SYNOPSYS_UNCONNECTED__154, 
        SYNOPSYS_UNCONNECTED__155, SYNOPSYS_UNCONNECTED__156, 
        SYNOPSYS_UNCONNECTED__157, SYNOPSYS_UNCONNECTED__158, 
        SYNOPSYS_UNCONNECTED__159, \add_out_s2[5][31] , \add_out_s2[5][30] , 
        \add_out_s2[5][29] , \add_out_s2[5][28] , \add_out_s2[5][27] , 
        \add_out_s2[5][26] , \add_out_s2[5][25] , \add_out_s2[5][24] , 
        \add_out_s2[5][23] , \add_out_s2[5][22] , \add_out_s2[5][21] , n13, 
        \add_out_s2[5][19] , \add_out_s2[5][18] , \add_out_s2[5][17] , 
        \add_out_s2[5][16] , \add_out_s2[5][15] , \add_out_s2[5][14] , 
        \add_out_s2[5][13] , \add_out_s2[5][12] , \add_out_s2[5][11] , 
        \add_out_s2[5][10] , \add_out_s2[5][9] , \add_out_s2[5][8] , 
        \add_out_s2[5][7] , \add_out_s2[5][6] , \add_out_s2[5][5] , 
        \add_out_s2[5][4] , \add_out_s2[5][3] , \add_out_s2[5][2] , 
        \add_out_s2[5][1] , \add_out_s2[5][0] }) );
  ADDER_P4_N_BIT64_10 adder_6 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, \mux_out[6][31] , \mux_out[6][30] , \mux_out[6][29] , 
        \mux_out[6][28] , \mux_out[6][27] , \mux_out[6][26] , \mux_out[6][25] , 
        \mux_out[6][24] , \mux_out[6][23] , \mux_out[6][22] , \mux_out[6][21] , 
        \mux_out[6][20] , \mux_out[6][19] , \mux_out[6][18] , \mux_out[6][17] , 
        \mux_out[6][16] , \mux_out[6][15] , \mux_out[6][14] , \mux_out[6][13] , 
        \mux_out[6][12] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        \add_out_s2[5][31] , \add_out_s2[5][30] , \add_out_s2[5][29] , 
        \add_out_s2[5][28] , \add_out_s2[5][27] , \add_out_s2[5][26] , 
        \add_out_s2[5][25] , \add_out_s2[5][24] , \add_out_s2[5][23] , 
        \add_out_s2[5][22] , \add_out_s2[5][21] , n13, \add_out_s2[5][19] , 
        \add_out_s2[5][18] , \add_out_s2[5][17] , \add_out_s2[5][16] , 
        \add_out_s2[5][15] , \add_out_s2[5][14] , \add_out_s2[5][13] , 
        \add_out_s2[5][12] , \add_out_s2[5][11] , \add_out_s2[5][10] , 
        \add_out_s2[5][9] , \add_out_s2[5][8] , \add_out_s2[5][7] , 
        \add_out_s2[5][6] , \add_out_s2[5][5] , \add_out_s2[5][4] , 
        \add_out_s2[5][3] , \add_out_s2[5][2] , \add_out_s2[5][1] , 
        \add_out_s2[5][0] }), .add_sub(1'b0), .SUM({SYNOPSYS_UNCONNECTED__160, 
        SYNOPSYS_UNCONNECTED__161, SYNOPSYS_UNCONNECTED__162, 
        SYNOPSYS_UNCONNECTED__163, SYNOPSYS_UNCONNECTED__164, 
        SYNOPSYS_UNCONNECTED__165, SYNOPSYS_UNCONNECTED__166, 
        SYNOPSYS_UNCONNECTED__167, SYNOPSYS_UNCONNECTED__168, 
        SYNOPSYS_UNCONNECTED__169, SYNOPSYS_UNCONNECTED__170, 
        SYNOPSYS_UNCONNECTED__171, SYNOPSYS_UNCONNECTED__172, 
        SYNOPSYS_UNCONNECTED__173, SYNOPSYS_UNCONNECTED__174, 
        SYNOPSYS_UNCONNECTED__175, SYNOPSYS_UNCONNECTED__176, 
        SYNOPSYS_UNCONNECTED__177, SYNOPSYS_UNCONNECTED__178, 
        SYNOPSYS_UNCONNECTED__179, SYNOPSYS_UNCONNECTED__180, 
        SYNOPSYS_UNCONNECTED__181, SYNOPSYS_UNCONNECTED__182, 
        SYNOPSYS_UNCONNECTED__183, SYNOPSYS_UNCONNECTED__184, 
        SYNOPSYS_UNCONNECTED__185, SYNOPSYS_UNCONNECTED__186, 
        SYNOPSYS_UNCONNECTED__187, SYNOPSYS_UNCONNECTED__188, 
        SYNOPSYS_UNCONNECTED__189, SYNOPSYS_UNCONNECTED__190, 
        SYNOPSYS_UNCONNECTED__191, \add_out_s2[6][31] , \add_out_s2[6][30] , 
        \add_out_s2[6][29] , \add_out_s2[6][28] , \add_out_s2[6][27] , 
        \add_out_s2[6][26] , \add_out_s2[6][25] , \add_out_s2[6][24] , 
        \add_out_s2[6][23] , \add_out_s2[6][22] , \add_out_s2[6][21] , 
        \add_out_s2[6][20] , \add_out_s2[6][19] , \add_out_s2[6][18] , 
        \add_out_s2[6][17] , \add_out_s2[6][16] , \add_out_s2[6][15] , 
        \add_out_s2[6][14] , \add_out_s2[6][13] , \add_out_s2[6][12] , 
        \add_out_s2[6][11] , \add_out_s2[6][10] , \add_out_s2[6][9] , 
        \add_out_s2[6][8] , \add_out_s2[6][7] , \add_out_s2[6][6] , 
        \add_out_s2[6][5] , \add_out_s2[6][4] , \add_out_s2[6][3] , 
        \add_out_s2[6][2] , \add_out_s2[6][1] , \add_out_s2[6][0] }) );
  ADDER_P4_N_BIT64_9 adder_7 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, \mux_out[7][31] , \mux_out[7][30] , \mux_out[7][29] , 
        \mux_out[7][28] , \mux_out[7][27] , \mux_out[7][26] , \mux_out[7][25] , 
        \mux_out[7][24] , \mux_out[7][23] , \mux_out[7][22] , \mux_out[7][21] , 
        \mux_out[7][20] , \mux_out[7][19] , \mux_out[7][18] , \mux_out[7][17] , 
        \mux_out[7][16] , \mux_out[7][15] , \mux_out[7][14] , 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        \add_out_s2[6][31] , \add_out_s2[6][30] , \add_out_s2[6][29] , 
        \add_out_s2[6][28] , \add_out_s2[6][27] , \add_out_s2[6][26] , 
        \add_out_s2[6][25] , \add_out_s2[6][24] , \add_out_s2[6][23] , 
        \add_out_s2[6][22] , \add_out_s2[6][21] , \add_out_s2[6][20] , 
        \add_out_s2[6][19] , \add_out_s2[6][18] , \add_out_s2[6][17] , 
        \add_out_s2[6][16] , \add_out_s2[6][15] , \add_out_s2[6][14] , 
        \add_out_s2[6][13] , \add_out_s2[6][12] , \add_out_s2[6][11] , 
        \add_out_s2[6][10] , \add_out_s2[6][9] , \add_out_s2[6][8] , 
        \add_out_s2[6][7] , \add_out_s2[6][6] , \add_out_s2[6][5] , 
        \add_out_s2[6][4] , \add_out_s2[6][3] , \add_out_s2[6][2] , 
        \add_out_s2[6][1] , \add_out_s2[6][0] }), .add_sub(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__192, SYNOPSYS_UNCONNECTED__193, 
        SYNOPSYS_UNCONNECTED__194, SYNOPSYS_UNCONNECTED__195, 
        SYNOPSYS_UNCONNECTED__196, SYNOPSYS_UNCONNECTED__197, 
        SYNOPSYS_UNCONNECTED__198, SYNOPSYS_UNCONNECTED__199, 
        SYNOPSYS_UNCONNECTED__200, SYNOPSYS_UNCONNECTED__201, 
        SYNOPSYS_UNCONNECTED__202, SYNOPSYS_UNCONNECTED__203, 
        SYNOPSYS_UNCONNECTED__204, SYNOPSYS_UNCONNECTED__205, 
        SYNOPSYS_UNCONNECTED__206, SYNOPSYS_UNCONNECTED__207, 
        SYNOPSYS_UNCONNECTED__208, SYNOPSYS_UNCONNECTED__209, 
        SYNOPSYS_UNCONNECTED__210, SYNOPSYS_UNCONNECTED__211, 
        SYNOPSYS_UNCONNECTED__212, SYNOPSYS_UNCONNECTED__213, 
        SYNOPSYS_UNCONNECTED__214, SYNOPSYS_UNCONNECTED__215, 
        SYNOPSYS_UNCONNECTED__216, SYNOPSYS_UNCONNECTED__217, 
        SYNOPSYS_UNCONNECTED__218, SYNOPSYS_UNCONNECTED__219, 
        SYNOPSYS_UNCONNECTED__220, SYNOPSYS_UNCONNECTED__221, 
        SYNOPSYS_UNCONNECTED__222, SYNOPSYS_UNCONNECTED__223, 
        \add_out_s2[7][31] , \add_out_s2[7][30] , \add_out_s2[7][29] , n14, 
        \add_out_s2[7][27] , \add_out_s2[7][26] , \add_out_s2[7][25] , 
        \add_out_s2[7][24] , \add_out_s2[7][23] , \add_out_s2[7][22] , 
        \add_out_s2[7][21] , \add_out_s2[7][20] , \add_out_s2[7][19] , 
        \add_out_s2[7][18] , \add_out_s2[7][17] , \add_out_s2[7][16] , 
        \add_out_s2[7][15] , \add_out_s2[7][14] , \add_out_s2[7][13] , 
        \add_out_s2[7][12] , \add_out_s2[7][11] , \add_out_s2[7][10] , 
        \add_out_s2[7][9] , \add_out_s2[7][8] , \add_out_s2[7][7] , 
        \add_out_s2[7][6] , \add_out_s2[7][5] , \add_out_s2[7][4] , 
        \add_out_s2[7][3] , \add_out_s2[7][2] , \add_out_s2[7][1] , 
        \add_out_s2[7][0] }) );
  ADDER_P4_N_BIT64_8 adder_8 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, \mux_out[8][31] , \mux_out[8][30] , \mux_out[8][29] , 
        \mux_out[8][28] , \mux_out[8][27] , \mux_out[8][26] , \mux_out[8][25] , 
        \mux_out[8][24] , \mux_out[8][23] , \mux_out[8][22] , \mux_out[8][21] , 
        \mux_out[8][20] , \mux_out[8][19] , \mux_out[8][18] , \mux_out[8][17] , 
        \mux_out[8][16] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, \add_out_s2[7][31] , \add_out_s2[7][30] , 
        \add_out_s2[7][29] , n14, \add_out_s2[7][27] , \add_out_s2[7][26] , 
        \add_out_s2[7][25] , \add_out_s2[7][24] , \add_out_s2[7][23] , 
        \add_out_s2[7][22] , \add_out_s2[7][21] , \add_out_s2[7][20] , 
        \add_out_s2[7][19] , \add_out_s2[7][18] , \add_out_s2[7][17] , 
        \add_out_s2[7][16] , \add_out_s2[7][15] , \add_out_s2[7][14] , 
        \add_out_s2[7][13] , \add_out_s2[7][12] , \add_out_s2[7][11] , 
        \add_out_s2[7][10] , \add_out_s2[7][9] , \add_out_s2[7][8] , 
        \add_out_s2[7][7] , \add_out_s2[7][6] , \add_out_s2[7][5] , 
        \add_out_s2[7][4] , \add_out_s2[7][3] , \add_out_s2[7][2] , 
        \add_out_s2[7][1] , \add_out_s2[7][0] }), .add_sub(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__224, SYNOPSYS_UNCONNECTED__225, 
        SYNOPSYS_UNCONNECTED__226, SYNOPSYS_UNCONNECTED__227, 
        SYNOPSYS_UNCONNECTED__228, SYNOPSYS_UNCONNECTED__229, 
        SYNOPSYS_UNCONNECTED__230, SYNOPSYS_UNCONNECTED__231, 
        SYNOPSYS_UNCONNECTED__232, SYNOPSYS_UNCONNECTED__233, 
        SYNOPSYS_UNCONNECTED__234, SYNOPSYS_UNCONNECTED__235, 
        SYNOPSYS_UNCONNECTED__236, SYNOPSYS_UNCONNECTED__237, 
        SYNOPSYS_UNCONNECTED__238, SYNOPSYS_UNCONNECTED__239, 
        SYNOPSYS_UNCONNECTED__240, SYNOPSYS_UNCONNECTED__241, 
        SYNOPSYS_UNCONNECTED__242, SYNOPSYS_UNCONNECTED__243, 
        SYNOPSYS_UNCONNECTED__244, SYNOPSYS_UNCONNECTED__245, 
        SYNOPSYS_UNCONNECTED__246, SYNOPSYS_UNCONNECTED__247, 
        SYNOPSYS_UNCONNECTED__248, SYNOPSYS_UNCONNECTED__249, 
        SYNOPSYS_UNCONNECTED__250, SYNOPSYS_UNCONNECTED__251, 
        SYNOPSYS_UNCONNECTED__252, SYNOPSYS_UNCONNECTED__253, 
        SYNOPSYS_UNCONNECTED__254, SYNOPSYS_UNCONNECTED__255, 
        \add_out_s2[8][31] , \add_out_s2[8][30] , \add_out_s2[8][29] , 
        \add_out_s2[8][28] , \add_out_s2[8][27] , \add_out_s2[8][26] , 
        \add_out_s2[8][25] , \add_out_s2[8][24] , \add_out_s2[8][23] , 
        \add_out_s2[8][22] , \add_out_s2[8][21] , \add_out_s2[8][20] , 
        \add_out_s2[8][19] , \add_out_s2[8][18] , \add_out_s2[8][17] , 
        \add_out_s2[8][16] , \add_out_s2[8][15] , \add_out_s2[8][14] , 
        \add_out_s2[8][13] , \add_out_s2[8][12] , \add_out_s2[8][11] , 
        \add_out_s2[8][10] , \add_out_s2[8][9] , \add_out_s2[8][8] , 
        \add_out_s2[8][7] , \add_out_s2[8][6] , \add_out_s2[8][5] , 
        \add_out_s2[8][4] , \add_out_s2[8][3] , \add_out_s2[8][2] , 
        \add_out_s2[8][1] , \add_out_s2[8][0] }) );
  ADDER_P4_N_BIT64_7 adder_9 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, \mux_out[9][31] , \mux_out[9][30] , \mux_out[9][29] , 
        \mux_out[9][28] , \mux_out[9][27] , \mux_out[9][26] , \mux_out[9][25] , 
        \mux_out[9][24] , \mux_out[9][23] , \mux_out[9][22] , \mux_out[9][21] , 
        \mux_out[9][20] , \mux_out[9][19] , \mux_out[9][18] , 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        \add_out_s3[8][31] , \add_out_s3[8][30] , \add_out_s3[8][29] , 
        \add_out_s3[8][28] , \add_out_s3[8][27] , \add_out_s3[8][26] , 
        \add_out_s3[8][25] , \add_out_s3[8][24] , \add_out_s3[8][23] , 
        \add_out_s3[8][22] , \add_out_s3[8][21] , \add_out_s3[8][20] , 
        \add_out_s3[8][19] , \add_out_s3[8][18] , \add_out_s3[8][17] , 
        \add_out_s3[8][16] , \add_out_s3[8][15] , \add_out_s3[8][14] , 
        \add_out_s3[8][13] , \add_out_s3[8][12] , \add_out_s3[8][11] , 
        \add_out_s3[8][10] , \add_out_s3[8][9] , \add_out_s3[8][8] , 
        \add_out_s3[8][7] , \add_out_s3[8][6] , \add_out_s3[8][5] , 
        \add_out_s3[8][4] , \add_out_s3[8][3] , \add_out_s3[8][2] , 
        \add_out_s3[8][1] , \add_out_s3[8][0] }), .add_sub(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__256, SYNOPSYS_UNCONNECTED__257, 
        SYNOPSYS_UNCONNECTED__258, SYNOPSYS_UNCONNECTED__259, 
        SYNOPSYS_UNCONNECTED__260, SYNOPSYS_UNCONNECTED__261, 
        SYNOPSYS_UNCONNECTED__262, SYNOPSYS_UNCONNECTED__263, 
        SYNOPSYS_UNCONNECTED__264, SYNOPSYS_UNCONNECTED__265, 
        SYNOPSYS_UNCONNECTED__266, SYNOPSYS_UNCONNECTED__267, 
        SYNOPSYS_UNCONNECTED__268, SYNOPSYS_UNCONNECTED__269, 
        SYNOPSYS_UNCONNECTED__270, SYNOPSYS_UNCONNECTED__271, 
        SYNOPSYS_UNCONNECTED__272, SYNOPSYS_UNCONNECTED__273, 
        SYNOPSYS_UNCONNECTED__274, SYNOPSYS_UNCONNECTED__275, 
        SYNOPSYS_UNCONNECTED__276, SYNOPSYS_UNCONNECTED__277, 
        SYNOPSYS_UNCONNECTED__278, SYNOPSYS_UNCONNECTED__279, 
        SYNOPSYS_UNCONNECTED__280, SYNOPSYS_UNCONNECTED__281, 
        SYNOPSYS_UNCONNECTED__282, SYNOPSYS_UNCONNECTED__283, 
        SYNOPSYS_UNCONNECTED__284, SYNOPSYS_UNCONNECTED__285, 
        SYNOPSYS_UNCONNECTED__286, SYNOPSYS_UNCONNECTED__287, 
        \add_out_s3[9][31] , \add_out_s3[9][30] , \add_out_s3[9][29] , 
        \add_out_s3[9][28] , \add_out_s3[9][27] , \add_out_s3[9][26] , 
        \add_out_s3[9][25] , \add_out_s3[9][24] , \add_out_s3[9][23] , 
        \add_out_s3[9][22] , \add_out_s3[9][21] , \add_out_s3[9][20] , 
        \add_out_s3[9][19] , \add_out_s3[9][18] , \add_out_s3[9][17] , 
        \add_out_s3[9][16] , \add_out_s3[9][15] , \add_out_s3[9][14] , 
        \add_out_s3[9][13] , \add_out_s3[9][12] , \add_out_s3[9][11] , 
        \add_out_s3[9][10] , \add_out_s3[9][9] , \add_out_s3[9][8] , 
        \add_out_s3[9][7] , \add_out_s3[9][6] , \add_out_s3[9][5] , 
        \add_out_s3[9][4] , \add_out_s3[9][3] , \add_out_s3[9][2] , 
        \add_out_s3[9][1] , \add_out_s3[9][0] }) );
  ADDER_P4_N_BIT64_6 adder_10 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, \mux_out[10][31] , \mux_out[10][30] , \mux_out[10][29] , 
        \mux_out[10][28] , \mux_out[10][27] , \mux_out[10][26] , 
        \mux_out[10][25] , \mux_out[10][24] , \mux_out[10][23] , 
        \mux_out[10][22] , \mux_out[10][21] , \mux_out[10][20] , 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, \add_out_s3[9][31] , \add_out_s3[9][30] , 
        \add_out_s3[9][29] , \add_out_s3[9][28] , \add_out_s3[9][27] , 
        \add_out_s3[9][26] , \add_out_s3[9][25] , \add_out_s3[9][24] , 
        \add_out_s3[9][23] , \add_out_s3[9][22] , \add_out_s3[9][21] , 
        \add_out_s3[9][20] , \add_out_s3[9][19] , \add_out_s3[9][18] , 
        \add_out_s3[9][17] , \add_out_s3[9][16] , \add_out_s3[9][15] , 
        \add_out_s3[9][14] , \add_out_s3[9][13] , \add_out_s3[9][12] , 
        \add_out_s3[9][11] , \add_out_s3[9][10] , \add_out_s3[9][9] , 
        \add_out_s3[9][8] , \add_out_s3[9][7] , \add_out_s3[9][6] , 
        \add_out_s3[9][5] , \add_out_s3[9][4] , \add_out_s3[9][3] , 
        \add_out_s3[9][2] , \add_out_s3[9][1] , \add_out_s3[9][0] }), 
        .add_sub(1'b0), .SUM({SYNOPSYS_UNCONNECTED__288, 
        SYNOPSYS_UNCONNECTED__289, SYNOPSYS_UNCONNECTED__290, 
        SYNOPSYS_UNCONNECTED__291, SYNOPSYS_UNCONNECTED__292, 
        SYNOPSYS_UNCONNECTED__293, SYNOPSYS_UNCONNECTED__294, 
        SYNOPSYS_UNCONNECTED__295, SYNOPSYS_UNCONNECTED__296, 
        SYNOPSYS_UNCONNECTED__297, SYNOPSYS_UNCONNECTED__298, 
        SYNOPSYS_UNCONNECTED__299, SYNOPSYS_UNCONNECTED__300, 
        SYNOPSYS_UNCONNECTED__301, SYNOPSYS_UNCONNECTED__302, 
        SYNOPSYS_UNCONNECTED__303, SYNOPSYS_UNCONNECTED__304, 
        SYNOPSYS_UNCONNECTED__305, SYNOPSYS_UNCONNECTED__306, 
        SYNOPSYS_UNCONNECTED__307, SYNOPSYS_UNCONNECTED__308, 
        SYNOPSYS_UNCONNECTED__309, SYNOPSYS_UNCONNECTED__310, 
        SYNOPSYS_UNCONNECTED__311, SYNOPSYS_UNCONNECTED__312, 
        SYNOPSYS_UNCONNECTED__313, SYNOPSYS_UNCONNECTED__314, 
        SYNOPSYS_UNCONNECTED__315, SYNOPSYS_UNCONNECTED__316, 
        SYNOPSYS_UNCONNECTED__317, SYNOPSYS_UNCONNECTED__318, 
        SYNOPSYS_UNCONNECTED__319, \add_out_s3[10][31] , \add_out_s3[10][30] , 
        \add_out_s3[10][29] , \add_out_s3[10][28] , \add_out_s3[10][27] , 
        \add_out_s3[10][26] , \add_out_s3[10][25] , \add_out_s3[10][24] , 
        \add_out_s3[10][23] , \add_out_s3[10][22] , \add_out_s3[10][21] , 
        \add_out_s3[10][20] , \add_out_s3[10][19] , \add_out_s3[10][18] , 
        \add_out_s3[10][17] , \add_out_s3[10][16] , \add_out_s3[10][15] , 
        \add_out_s3[10][14] , \add_out_s3[10][13] , \add_out_s3[10][12] , 
        \add_out_s3[10][11] , \add_out_s3[10][10] , \add_out_s3[10][9] , 
        \add_out_s3[10][8] , \add_out_s3[10][7] , \add_out_s3[10][6] , 
        \add_out_s3[10][5] , \add_out_s3[10][4] , \add_out_s3[10][3] , 
        \add_out_s3[10][2] , \add_out_s3[10][1] , \add_out_s3[10][0] }) );
  ADDER_P4_N_BIT64_5 adder_11 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, \mux_out[11][31] , \mux_out[11][30] , \mux_out[11][29] , 
        \mux_out[11][28] , \mux_out[11][27] , \mux_out[11][26] , 
        \mux_out[11][25] , \mux_out[11][24] , \mux_out[11][23] , 
        \mux_out[11][22] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        \add_out_s3[10][31] , \add_out_s3[10][30] , \add_out_s3[10][29] , 
        \add_out_s3[10][28] , \add_out_s3[10][27] , \add_out_s3[10][26] , 
        \add_out_s3[10][25] , \add_out_s3[10][24] , \add_out_s3[10][23] , 
        \add_out_s3[10][22] , \add_out_s3[10][21] , \add_out_s3[10][20] , 
        \add_out_s3[10][19] , \add_out_s3[10][18] , \add_out_s3[10][17] , 
        \add_out_s3[10][16] , \add_out_s3[10][15] , \add_out_s3[10][14] , 
        \add_out_s3[10][13] , \add_out_s3[10][12] , \add_out_s3[10][11] , 
        \add_out_s3[10][10] , \add_out_s3[10][9] , \add_out_s3[10][8] , 
        \add_out_s3[10][7] , \add_out_s3[10][6] , \add_out_s3[10][5] , 
        \add_out_s3[10][4] , \add_out_s3[10][3] , \add_out_s3[10][2] , 
        \add_out_s3[10][1] , \add_out_s3[10][0] }), .add_sub(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__320, SYNOPSYS_UNCONNECTED__321, 
        SYNOPSYS_UNCONNECTED__322, SYNOPSYS_UNCONNECTED__323, 
        SYNOPSYS_UNCONNECTED__324, SYNOPSYS_UNCONNECTED__325, 
        SYNOPSYS_UNCONNECTED__326, SYNOPSYS_UNCONNECTED__327, 
        SYNOPSYS_UNCONNECTED__328, SYNOPSYS_UNCONNECTED__329, 
        SYNOPSYS_UNCONNECTED__330, SYNOPSYS_UNCONNECTED__331, 
        SYNOPSYS_UNCONNECTED__332, SYNOPSYS_UNCONNECTED__333, 
        SYNOPSYS_UNCONNECTED__334, SYNOPSYS_UNCONNECTED__335, 
        SYNOPSYS_UNCONNECTED__336, SYNOPSYS_UNCONNECTED__337, 
        SYNOPSYS_UNCONNECTED__338, SYNOPSYS_UNCONNECTED__339, 
        SYNOPSYS_UNCONNECTED__340, SYNOPSYS_UNCONNECTED__341, 
        SYNOPSYS_UNCONNECTED__342, SYNOPSYS_UNCONNECTED__343, 
        SYNOPSYS_UNCONNECTED__344, SYNOPSYS_UNCONNECTED__345, 
        SYNOPSYS_UNCONNECTED__346, SYNOPSYS_UNCONNECTED__347, 
        SYNOPSYS_UNCONNECTED__348, SYNOPSYS_UNCONNECTED__349, 
        SYNOPSYS_UNCONNECTED__350, SYNOPSYS_UNCONNECTED__351, 
        \add_out_s3[11][31] , \add_out_s3[11][30] , \add_out_s3[11][29] , 
        \add_out_s3[11][28] , \add_out_s3[11][27] , \add_out_s3[11][26] , 
        \add_out_s3[11][25] , \add_out_s3[11][24] , \add_out_s3[11][23] , 
        \add_out_s3[11][22] , \add_out_s3[11][21] , \add_out_s3[11][20] , 
        \add_out_s3[11][19] , \add_out_s3[11][18] , \add_out_s3[11][17] , 
        \add_out_s3[11][16] , \add_out_s3[11][15] , \add_out_s3[11][14] , 
        \add_out_s3[11][13] , \add_out_s3[11][12] , \add_out_s3[11][11] , 
        \add_out_s3[11][10] , \add_out_s3[11][9] , \add_out_s3[11][8] , 
        \add_out_s3[11][7] , \add_out_s3[11][6] , \add_out_s3[11][5] , 
        \add_out_s3[11][4] , \add_out_s3[11][3] , \add_out_s3[11][2] , 
        \add_out_s3[11][1] , \add_out_s3[11][0] }) );
  ADDER_P4_N_BIT64_4 adder_12 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, \mux_out[12][31] , \mux_out[12][30] , \mux_out[12][29] , 
        \mux_out[12][28] , \mux_out[12][27] , \mux_out[12][26] , 
        \mux_out[12][25] , \mux_out[12][24] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, \add_out_s3[11][31] , \add_out_s3[11][30] , 
        \add_out_s3[11][29] , \add_out_s3[11][28] , \add_out_s3[11][27] , 
        \add_out_s3[11][26] , \add_out_s3[11][25] , \add_out_s3[11][24] , 
        \add_out_s3[11][23] , \add_out_s3[11][22] , \add_out_s3[11][21] , 
        \add_out_s3[11][20] , \add_out_s3[11][19] , \add_out_s3[11][18] , 
        \add_out_s3[11][17] , \add_out_s3[11][16] , \add_out_s3[11][15] , 
        \add_out_s3[11][14] , \add_out_s3[11][13] , \add_out_s3[11][12] , 
        \add_out_s3[11][11] , \add_out_s3[11][10] , \add_out_s3[11][9] , 
        \add_out_s3[11][8] , \add_out_s3[11][7] , \add_out_s3[11][6] , 
        \add_out_s3[11][5] , \add_out_s3[11][4] , \add_out_s3[11][3] , 
        \add_out_s3[11][2] , \add_out_s3[11][1] , \add_out_s3[11][0] }), 
        .add_sub(1'b0), .SUM({SYNOPSYS_UNCONNECTED__352, 
        SYNOPSYS_UNCONNECTED__353, SYNOPSYS_UNCONNECTED__354, 
        SYNOPSYS_UNCONNECTED__355, SYNOPSYS_UNCONNECTED__356, 
        SYNOPSYS_UNCONNECTED__357, SYNOPSYS_UNCONNECTED__358, 
        SYNOPSYS_UNCONNECTED__359, SYNOPSYS_UNCONNECTED__360, 
        SYNOPSYS_UNCONNECTED__361, SYNOPSYS_UNCONNECTED__362, 
        SYNOPSYS_UNCONNECTED__363, SYNOPSYS_UNCONNECTED__364, 
        SYNOPSYS_UNCONNECTED__365, SYNOPSYS_UNCONNECTED__366, 
        SYNOPSYS_UNCONNECTED__367, SYNOPSYS_UNCONNECTED__368, 
        SYNOPSYS_UNCONNECTED__369, SYNOPSYS_UNCONNECTED__370, 
        SYNOPSYS_UNCONNECTED__371, SYNOPSYS_UNCONNECTED__372, 
        SYNOPSYS_UNCONNECTED__373, SYNOPSYS_UNCONNECTED__374, 
        SYNOPSYS_UNCONNECTED__375, SYNOPSYS_UNCONNECTED__376, 
        SYNOPSYS_UNCONNECTED__377, SYNOPSYS_UNCONNECTED__378, 
        SYNOPSYS_UNCONNECTED__379, SYNOPSYS_UNCONNECTED__380, 
        SYNOPSYS_UNCONNECTED__381, SYNOPSYS_UNCONNECTED__382, 
        SYNOPSYS_UNCONNECTED__383, \add_out_s3[12][31] , \add_out_s3[12][30] , 
        \add_out_s3[12][29] , \add_out_s3[12][28] , \add_out_s3[12][27] , 
        \add_out_s3[12][26] , \add_out_s3[12][25] , \add_out_s3[12][24] , 
        \add_out_s3[12][23] , \add_out_s3[12][22] , \add_out_s3[12][21] , 
        \add_out_s3[12][20] , \add_out_s3[12][19] , \add_out_s3[12][18] , 
        \add_out_s3[12][17] , \add_out_s3[12][16] , \add_out_s3[12][15] , 
        \add_out_s3[12][14] , \add_out_s3[12][13] , \add_out_s3[12][12] , 
        \add_out_s3[12][11] , \add_out_s3[12][10] , \add_out_s3[12][9] , 
        \add_out_s3[12][8] , \add_out_s3[12][7] , \add_out_s3[12][6] , 
        \add_out_s3[12][5] , \add_out_s3[12][4] , \add_out_s3[12][3] , 
        \add_out_s3[12][2] , \add_out_s3[12][1] , \add_out_s3[12][0] }) );
  ADDER_P4_N_BIT64_3 adder_13 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, \mux_out[13][31] , \mux_out[13][30] , \mux_out[13][29] , 
        \mux_out[13][28] , \mux_out[13][27] , \mux_out[13][26] , 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \add_out_s4[12][31] , 
        \add_out_s4[12][30] , \add_out_s4[12][29] , \add_out_s4[12][28] , 
        \add_out_s4[12][27] , \add_out_s4[12][26] , \add_out_s4[12][25] , 
        \add_out_s4[12][24] , \add_out_s4[12][23] , \add_out_s4[12][22] , 
        \add_out_s4[12][21] , \add_out_s4[12][20] , \add_out_s4[12][19] , 
        \add_out_s4[12][18] , \add_out_s4[12][17] , \add_out_s4[12][16] , 
        \add_out_s4[12][15] , \add_out_s4[12][14] , \add_out_s4[12][13] , 
        \add_out_s4[12][12] , \add_out_s4[12][11] , \add_out_s4[12][10] , 
        \add_out_s4[12][9] , \add_out_s4[12][8] , \add_out_s4[12][7] , 
        \add_out_s4[12][6] , \add_out_s4[12][5] , \add_out_s4[12][4] , 
        \add_out_s4[12][3] , \add_out_s4[12][2] , \add_out_s4[12][1] , 
        \add_out_s4[12][0] }), .add_sub(1'b0), .SUM({SYNOPSYS_UNCONNECTED__384, 
        SYNOPSYS_UNCONNECTED__385, SYNOPSYS_UNCONNECTED__386, 
        SYNOPSYS_UNCONNECTED__387, SYNOPSYS_UNCONNECTED__388, 
        SYNOPSYS_UNCONNECTED__389, SYNOPSYS_UNCONNECTED__390, 
        SYNOPSYS_UNCONNECTED__391, SYNOPSYS_UNCONNECTED__392, 
        SYNOPSYS_UNCONNECTED__393, SYNOPSYS_UNCONNECTED__394, 
        SYNOPSYS_UNCONNECTED__395, SYNOPSYS_UNCONNECTED__396, 
        SYNOPSYS_UNCONNECTED__397, SYNOPSYS_UNCONNECTED__398, 
        SYNOPSYS_UNCONNECTED__399, SYNOPSYS_UNCONNECTED__400, 
        SYNOPSYS_UNCONNECTED__401, SYNOPSYS_UNCONNECTED__402, 
        SYNOPSYS_UNCONNECTED__403, SYNOPSYS_UNCONNECTED__404, 
        SYNOPSYS_UNCONNECTED__405, SYNOPSYS_UNCONNECTED__406, 
        SYNOPSYS_UNCONNECTED__407, SYNOPSYS_UNCONNECTED__408, 
        SYNOPSYS_UNCONNECTED__409, SYNOPSYS_UNCONNECTED__410, 
        SYNOPSYS_UNCONNECTED__411, SYNOPSYS_UNCONNECTED__412, 
        SYNOPSYS_UNCONNECTED__413, SYNOPSYS_UNCONNECTED__414, 
        SYNOPSYS_UNCONNECTED__415, \add_out_s4[13][31] , \add_out_s4[13][30] , 
        \add_out_s4[13][29] , \add_out_s4[13][28] , \add_out_s4[13][27] , 
        \add_out_s4[13][26] , \add_out_s4[13][25] , \add_out_s4[13][24] , 
        \add_out_s4[13][23] , \add_out_s4[13][22] , \add_out_s4[13][21] , 
        \add_out_s4[13][20] , \add_out_s4[13][19] , \add_out_s4[13][18] , 
        \add_out_s4[13][17] , \add_out_s4[13][16] , \add_out_s4[13][15] , 
        \add_out_s4[13][14] , \add_out_s4[13][13] , \add_out_s4[13][12] , 
        \add_out_s4[13][11] , \add_out_s4[13][10] , \add_out_s4[13][9] , 
        \add_out_s4[13][8] , \add_out_s4[13][7] , \add_out_s4[13][6] , 
        \add_out_s4[13][5] , \add_out_s4[13][4] , \add_out_s4[13][3] , 
        \add_out_s4[13][2] , \add_out_s4[13][1] , \add_out_s4[13][0] }) );
  ADDER_P4_N_BIT64_2 adder_14 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, \mux_out[14][31] , \mux_out[14][30] , \mux_out[14][29] , 
        \mux_out[14][28] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \add_out_s4[13][31] , 
        \add_out_s4[13][30] , \add_out_s4[13][29] , \add_out_s4[13][28] , 
        \add_out_s4[13][27] , \add_out_s4[13][26] , \add_out_s4[13][25] , 
        \add_out_s4[13][24] , \add_out_s4[13][23] , \add_out_s4[13][22] , 
        \add_out_s4[13][21] , \add_out_s4[13][20] , \add_out_s4[13][19] , 
        \add_out_s4[13][18] , \add_out_s4[13][17] , \add_out_s4[13][16] , 
        \add_out_s4[13][15] , \add_out_s4[13][14] , \add_out_s4[13][13] , 
        \add_out_s4[13][12] , \add_out_s4[13][11] , \add_out_s4[13][10] , 
        \add_out_s4[13][9] , \add_out_s4[13][8] , \add_out_s4[13][7] , 
        \add_out_s4[13][6] , \add_out_s4[13][5] , \add_out_s4[13][4] , 
        \add_out_s4[13][3] , \add_out_s4[13][2] , \add_out_s4[13][1] , 
        \add_out_s4[13][0] }), .add_sub(1'b0), .SUM({SYNOPSYS_UNCONNECTED__416, 
        SYNOPSYS_UNCONNECTED__417, SYNOPSYS_UNCONNECTED__418, 
        SYNOPSYS_UNCONNECTED__419, SYNOPSYS_UNCONNECTED__420, 
        SYNOPSYS_UNCONNECTED__421, SYNOPSYS_UNCONNECTED__422, 
        SYNOPSYS_UNCONNECTED__423, SYNOPSYS_UNCONNECTED__424, 
        SYNOPSYS_UNCONNECTED__425, SYNOPSYS_UNCONNECTED__426, 
        SYNOPSYS_UNCONNECTED__427, SYNOPSYS_UNCONNECTED__428, 
        SYNOPSYS_UNCONNECTED__429, SYNOPSYS_UNCONNECTED__430, 
        SYNOPSYS_UNCONNECTED__431, SYNOPSYS_UNCONNECTED__432, 
        SYNOPSYS_UNCONNECTED__433, SYNOPSYS_UNCONNECTED__434, 
        SYNOPSYS_UNCONNECTED__435, SYNOPSYS_UNCONNECTED__436, 
        SYNOPSYS_UNCONNECTED__437, SYNOPSYS_UNCONNECTED__438, 
        SYNOPSYS_UNCONNECTED__439, SYNOPSYS_UNCONNECTED__440, 
        SYNOPSYS_UNCONNECTED__441, SYNOPSYS_UNCONNECTED__442, 
        SYNOPSYS_UNCONNECTED__443, SYNOPSYS_UNCONNECTED__444, 
        SYNOPSYS_UNCONNECTED__445, SYNOPSYS_UNCONNECTED__446, 
        SYNOPSYS_UNCONNECTED__447, \add_out_s4[14][31] , \add_out_s4[14][30] , 
        \add_out_s4[14][29] , \add_out_s4[14][28] , \add_out_s4[14][27] , 
        \add_out_s4[14][26] , \add_out_s4[14][25] , \add_out_s4[14][24] , 
        \add_out_s4[14][23] , \add_out_s4[14][22] , \add_out_s4[14][21] , 
        \add_out_s4[14][20] , \add_out_s4[14][19] , \add_out_s4[14][18] , 
        \add_out_s4[14][17] , \add_out_s4[14][16] , \add_out_s4[14][15] , 
        \add_out_s4[14][14] , \add_out_s4[14][13] , \add_out_s4[14][12] , 
        \add_out_s4[14][11] , \add_out_s4[14][10] , \add_out_s4[14][9] , 
        \add_out_s4[14][8] , \add_out_s4[14][7] , \add_out_s4[14][6] , 
        \add_out_s4[14][5] , \add_out_s4[14][4] , \add_out_s4[14][3] , 
        \add_out_s4[14][2] , \add_out_s4[14][1] , \add_out_s4[14][0] }) );
  ADDER_P4_N_BIT64_1 adder_15 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, \mux_out[15][31] , \mux_out[15][30] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        \add_out_s4[14][31] , \add_out_s4[14][30] , \add_out_s4[14][29] , 
        \add_out_s4[14][28] , \add_out_s4[14][27] , \add_out_s4[14][26] , 
        \add_out_s4[14][25] , \add_out_s4[14][24] , \add_out_s4[14][23] , 
        \add_out_s4[14][22] , \add_out_s4[14][21] , \add_out_s4[14][20] , 
        \add_out_s4[14][19] , \add_out_s4[14][18] , \add_out_s4[14][17] , 
        \add_out_s4[14][16] , \add_out_s4[14][15] , \add_out_s4[14][14] , 
        \add_out_s4[14][13] , \add_out_s4[14][12] , \add_out_s4[14][11] , 
        \add_out_s4[14][10] , \add_out_s4[14][9] , \add_out_s4[14][8] , 
        \add_out_s4[14][7] , \add_out_s4[14][6] , \add_out_s4[14][5] , 
        \add_out_s4[14][4] , \add_out_s4[14][3] , \add_out_s4[14][2] , 
        \add_out_s4[14][1] , \add_out_s4[14][0] }), .add_sub(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__448, SYNOPSYS_UNCONNECTED__449, 
        SYNOPSYS_UNCONNECTED__450, SYNOPSYS_UNCONNECTED__451, 
        SYNOPSYS_UNCONNECTED__452, SYNOPSYS_UNCONNECTED__453, 
        SYNOPSYS_UNCONNECTED__454, SYNOPSYS_UNCONNECTED__455, 
        SYNOPSYS_UNCONNECTED__456, SYNOPSYS_UNCONNECTED__457, 
        SYNOPSYS_UNCONNECTED__458, SYNOPSYS_UNCONNECTED__459, 
        SYNOPSYS_UNCONNECTED__460, SYNOPSYS_UNCONNECTED__461, 
        SYNOPSYS_UNCONNECTED__462, SYNOPSYS_UNCONNECTED__463, 
        SYNOPSYS_UNCONNECTED__464, SYNOPSYS_UNCONNECTED__465, 
        SYNOPSYS_UNCONNECTED__466, SYNOPSYS_UNCONNECTED__467, 
        SYNOPSYS_UNCONNECTED__468, SYNOPSYS_UNCONNECTED__469, 
        SYNOPSYS_UNCONNECTED__470, SYNOPSYS_UNCONNECTED__471, 
        SYNOPSYS_UNCONNECTED__472, SYNOPSYS_UNCONNECTED__473, 
        SYNOPSYS_UNCONNECTED__474, SYNOPSYS_UNCONNECTED__475, 
        SYNOPSYS_UNCONNECTED__476, SYNOPSYS_UNCONNECTED__477, 
        SYNOPSYS_UNCONNECTED__478, SYNOPSYS_UNCONNECTED__479, P[31:0]}) );
  MUX_8to1_N64_0 mux_0 ( .IN0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, A[31:24], \sub_x_1/B[23] , 
        \sub_x_1/B[22] , \sub_x_1/B[21] , A[20:18], \sub_x_1/B[17] , A[16], 
        \sub_x_1/B[15] , A[14:12], n643, n642, A[9], n641, n640, n639, n638, 
        n637, n626, n625, n636, n635}), .IN2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, \A_shifted[-32][62] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .IN3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN4({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \A_shifted[-32][61] , 
        \A_shifted[-32][60] , \A_shifted[-32][59] , \A_shifted[-32][58] , 
        \A_shifted[-32][57] , \A_shifted[-32][56] , \A_shifted[-32][55] , 
        \A_shifted[-32][54] , \A_shifted[-32][53] , \A_shifted[-32][52] , 
        \A_shifted[-32][51] , \A_shifted[-32][50] , \A_shifted[-32][49] , 
        \A_shifted[-32][48] , \A_shifted[-32][47] , \A_shifted[-32][46] , 
        \A_shifted[-32][45] , n91, \A_shifted[-32][43] , \A_shifted[-32][42] , 
        \A_shifted[-32][41] , \A_shifted[-32][40] , n634, n632, n17, n630, n19, 
        n23, n18, n628, 1'b0, 1'b0}), .IN5({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN6({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .IN7({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .SEL({
        \encoder_out[0][2] , \encoder_out[0][1] , \encoder_out[0][0] }), .Y({
        SYNOPSYS_UNCONNECTED__480, SYNOPSYS_UNCONNECTED__481, 
        SYNOPSYS_UNCONNECTED__482, SYNOPSYS_UNCONNECTED__483, 
        SYNOPSYS_UNCONNECTED__484, SYNOPSYS_UNCONNECTED__485, 
        SYNOPSYS_UNCONNECTED__486, SYNOPSYS_UNCONNECTED__487, 
        SYNOPSYS_UNCONNECTED__488, SYNOPSYS_UNCONNECTED__489, 
        SYNOPSYS_UNCONNECTED__490, SYNOPSYS_UNCONNECTED__491, 
        SYNOPSYS_UNCONNECTED__492, SYNOPSYS_UNCONNECTED__493, 
        SYNOPSYS_UNCONNECTED__494, SYNOPSYS_UNCONNECTED__495, 
        SYNOPSYS_UNCONNECTED__496, SYNOPSYS_UNCONNECTED__497, 
        SYNOPSYS_UNCONNECTED__498, SYNOPSYS_UNCONNECTED__499, 
        SYNOPSYS_UNCONNECTED__500, SYNOPSYS_UNCONNECTED__501, 
        SYNOPSYS_UNCONNECTED__502, SYNOPSYS_UNCONNECTED__503, 
        SYNOPSYS_UNCONNECTED__504, SYNOPSYS_UNCONNECTED__505, 
        SYNOPSYS_UNCONNECTED__506, SYNOPSYS_UNCONNECTED__507, 
        SYNOPSYS_UNCONNECTED__508, SYNOPSYS_UNCONNECTED__509, 
        SYNOPSYS_UNCONNECTED__510, SYNOPSYS_UNCONNECTED__511, 
        \add_out_s1[0][31] , \add_out_s1[0][30] , \add_out_s1[0][29] , 
        \add_out_s1[0][28] , \add_out_s1[0][27] , \add_out_s1[0][26] , 
        \add_out_s1[0][25] , \add_out_s1[0][24] , \add_out_s1[0][23] , 
        \add_out_s1[0][22] , \add_out_s1[0][21] , \add_out_s1[0][20] , 
        \add_out_s1[0][19] , \add_out_s1[0][18] , \add_out_s1[0][17] , 
        \add_out_s1[0][16] , \add_out_s1[0][15] , \add_out_s1[0][14] , 
        \add_out_s1[0][13] , \add_out_s1[0][12] , \add_out_s1[0][11] , 
        \add_out_s1[0][10] , \add_out_s1[0][9] , \add_out_s1[0][8] , 
        \add_out_s1[0][7] , \add_out_s1[0][6] , \add_out_s1[0][5] , 
        \add_out_s1[0][4] , \add_out_s1[0][3] , \add_out_s1[0][2] , 
        \add_out_s1[0][1] , \add_out_s1[0][0] }) );
  MUX_8to1_N64_15 mux_1 ( .IN0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, A[29:24], \sub_x_1/B[23] , 
        \sub_x_1/B[22] , \sub_x_1/B[21] , A[20:18], \sub_x_1/B[17] , A[16], 
        \sub_x_1/B[15] , A[14:12], n643, n642, A[9], n641, n640, n639, n638, 
        n637, n626, n625, n636, n635, 1'b0, 1'b0}), .IN2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \A_shifted[-32][60] , 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .IN3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN4({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \A_shifted[-32][59] , 
        n56, \A_shifted[-32][57] , \A_shifted[-32][56] , \A_shifted[-32][55] , 
        \A_shifted[-32][54] , \A_shifted[-32][53] , \A_shifted[-32][52] , 
        \A_shifted[-32][51] , \A_shifted[-32][50] , \A_shifted[-32][49] , 
        \A_shifted[-32][48] , \A_shifted[-32][47] , \A_shifted[-32][46] , 
        \A_shifted[-32][45] , n91, \A_shifted[-32][43] , \A_shifted[-32][42] , 
        \A_shifted[-32][41] , \A_shifted[-32][40] , n633, n631, n17, n629, n19, 
        n23, n18, n628, 1'b0, 1'b0, 1'b0, 1'b0}), .IN5({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN6({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN7({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL({\encoder_out[1][2] , \encoder_out[1][1] , \encoder_out[1][0] }), 
        .Y({SYNOPSYS_UNCONNECTED__512, SYNOPSYS_UNCONNECTED__513, 
        SYNOPSYS_UNCONNECTED__514, SYNOPSYS_UNCONNECTED__515, 
        SYNOPSYS_UNCONNECTED__516, SYNOPSYS_UNCONNECTED__517, 
        SYNOPSYS_UNCONNECTED__518, SYNOPSYS_UNCONNECTED__519, 
        SYNOPSYS_UNCONNECTED__520, SYNOPSYS_UNCONNECTED__521, 
        SYNOPSYS_UNCONNECTED__522, SYNOPSYS_UNCONNECTED__523, 
        SYNOPSYS_UNCONNECTED__524, SYNOPSYS_UNCONNECTED__525, 
        SYNOPSYS_UNCONNECTED__526, SYNOPSYS_UNCONNECTED__527, 
        SYNOPSYS_UNCONNECTED__528, SYNOPSYS_UNCONNECTED__529, 
        SYNOPSYS_UNCONNECTED__530, SYNOPSYS_UNCONNECTED__531, 
        SYNOPSYS_UNCONNECTED__532, SYNOPSYS_UNCONNECTED__533, 
        SYNOPSYS_UNCONNECTED__534, SYNOPSYS_UNCONNECTED__535, 
        SYNOPSYS_UNCONNECTED__536, SYNOPSYS_UNCONNECTED__537, 
        SYNOPSYS_UNCONNECTED__538, SYNOPSYS_UNCONNECTED__539, 
        SYNOPSYS_UNCONNECTED__540, SYNOPSYS_UNCONNECTED__541, 
        SYNOPSYS_UNCONNECTED__542, SYNOPSYS_UNCONNECTED__543, \mux_out[1][31] , 
        \mux_out[1][30] , \mux_out[1][29] , \mux_out[1][28] , \mux_out[1][27] , 
        \mux_out[1][26] , \mux_out[1][25] , \mux_out[1][24] , \mux_out[1][23] , 
        \mux_out[1][22] , \mux_out[1][21] , \mux_out[1][20] , \mux_out[1][19] , 
        \mux_out[1][18] , \mux_out[1][17] , \mux_out[1][16] , \mux_out[1][15] , 
        \mux_out[1][14] , \mux_out[1][13] , \mux_out[1][12] , \mux_out[1][11] , 
        \mux_out[1][10] , \mux_out[1][9] , \mux_out[1][8] , \mux_out[1][7] , 
        \mux_out[1][6] , \mux_out[1][5] , \mux_out[1][4] , \mux_out[1][3] , 
        \mux_out[1][2] , SYNOPSYS_UNCONNECTED__544, SYNOPSYS_UNCONNECTED__545}) );
  MUX_8to1_N64_14 mux_2 ( .IN0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, A[27:24], \sub_x_1/B[23] , 
        \sub_x_1/B[22] , \sub_x_1/B[21] , A[20:18], \sub_x_1/B[17] , A[16], 
        \sub_x_1/B[15] , A[14:12], n643, n642, A[9], n641, n640, n639, n638, 
        n637, n626, n625, n636, n635, 1'b0, 1'b0, 1'b0, 1'b0}), .IN2({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n56, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .IN3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN4({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \A_shifted[-32][57] , 
        \A_shifted[-32][56] , \A_shifted[-32][55] , n57, n32, n53, n33, n95, 
        n41, n93, n90, n50, n52, n92, n55, n96, n94, n54, n633, n631, n17, 
        n629, n19, n23, n18, n628, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN5(
        {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN6({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .IN7({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .SEL({\encoder_out[2][2] , 
        \encoder_out[2][1] , \encoder_out[2][0] }), .Y({
        SYNOPSYS_UNCONNECTED__546, SYNOPSYS_UNCONNECTED__547, 
        SYNOPSYS_UNCONNECTED__548, SYNOPSYS_UNCONNECTED__549, 
        SYNOPSYS_UNCONNECTED__550, SYNOPSYS_UNCONNECTED__551, 
        SYNOPSYS_UNCONNECTED__552, SYNOPSYS_UNCONNECTED__553, 
        SYNOPSYS_UNCONNECTED__554, SYNOPSYS_UNCONNECTED__555, 
        SYNOPSYS_UNCONNECTED__556, SYNOPSYS_UNCONNECTED__557, 
        SYNOPSYS_UNCONNECTED__558, SYNOPSYS_UNCONNECTED__559, 
        SYNOPSYS_UNCONNECTED__560, SYNOPSYS_UNCONNECTED__561, 
        SYNOPSYS_UNCONNECTED__562, SYNOPSYS_UNCONNECTED__563, 
        SYNOPSYS_UNCONNECTED__564, SYNOPSYS_UNCONNECTED__565, 
        SYNOPSYS_UNCONNECTED__566, SYNOPSYS_UNCONNECTED__567, 
        SYNOPSYS_UNCONNECTED__568, SYNOPSYS_UNCONNECTED__569, 
        SYNOPSYS_UNCONNECTED__570, SYNOPSYS_UNCONNECTED__571, 
        SYNOPSYS_UNCONNECTED__572, SYNOPSYS_UNCONNECTED__573, 
        SYNOPSYS_UNCONNECTED__574, SYNOPSYS_UNCONNECTED__575, 
        SYNOPSYS_UNCONNECTED__576, SYNOPSYS_UNCONNECTED__577, \mux_out[2][31] , 
        \mux_out[2][30] , \mux_out[2][29] , \mux_out[2][28] , \mux_out[2][27] , 
        \mux_out[2][26] , \mux_out[2][25] , \mux_out[2][24] , \mux_out[2][23] , 
        \mux_out[2][22] , \mux_out[2][21] , \mux_out[2][20] , \mux_out[2][19] , 
        \mux_out[2][18] , \mux_out[2][17] , \mux_out[2][16] , \mux_out[2][15] , 
        \mux_out[2][14] , \mux_out[2][13] , \mux_out[2][12] , \mux_out[2][11] , 
        \mux_out[2][10] , \mux_out[2][9] , \mux_out[2][8] , \mux_out[2][7] , 
        \mux_out[2][6] , \mux_out[2][5] , \mux_out[2][4] , 
        SYNOPSYS_UNCONNECTED__578, SYNOPSYS_UNCONNECTED__579, 
        SYNOPSYS_UNCONNECTED__580, SYNOPSYS_UNCONNECTED__581}) );
  MUX_8to1_N64_13 mux_3 ( .IN0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, A[25:24], \sub_x_1/B[23] , 
        \sub_x_1/B[22] , \sub_x_1/B[21] , A[20:18], \sub_x_1/B[17] , A[16], 
        \sub_x_1/B[15] , A[14:12], n643, n642, A[9], n641, n640, n639, n638, 
        n637, n626, n625, n636, n635, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .IN2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        \A_shifted[-32][56] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .IN3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN4({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, \A_shifted[-32][55] , n57, n32, n53, n33, n95, n41, 
        n93, n90, n50, n52, n92, n55, n96, n94, n54, n633, n631, n17, n630, 
        n19, n23, n18, n628, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .IN5({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN6({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .IN7({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .SEL({\encoder_out[3][2] , 
        \encoder_out[3][1] , \encoder_out[3][0] }), .Y({
        SYNOPSYS_UNCONNECTED__582, SYNOPSYS_UNCONNECTED__583, 
        SYNOPSYS_UNCONNECTED__584, SYNOPSYS_UNCONNECTED__585, 
        SYNOPSYS_UNCONNECTED__586, SYNOPSYS_UNCONNECTED__587, 
        SYNOPSYS_UNCONNECTED__588, SYNOPSYS_UNCONNECTED__589, 
        SYNOPSYS_UNCONNECTED__590, SYNOPSYS_UNCONNECTED__591, 
        SYNOPSYS_UNCONNECTED__592, SYNOPSYS_UNCONNECTED__593, 
        SYNOPSYS_UNCONNECTED__594, SYNOPSYS_UNCONNECTED__595, 
        SYNOPSYS_UNCONNECTED__596, SYNOPSYS_UNCONNECTED__597, 
        SYNOPSYS_UNCONNECTED__598, SYNOPSYS_UNCONNECTED__599, 
        SYNOPSYS_UNCONNECTED__600, SYNOPSYS_UNCONNECTED__601, 
        SYNOPSYS_UNCONNECTED__602, SYNOPSYS_UNCONNECTED__603, 
        SYNOPSYS_UNCONNECTED__604, SYNOPSYS_UNCONNECTED__605, 
        SYNOPSYS_UNCONNECTED__606, SYNOPSYS_UNCONNECTED__607, 
        SYNOPSYS_UNCONNECTED__608, SYNOPSYS_UNCONNECTED__609, 
        SYNOPSYS_UNCONNECTED__610, SYNOPSYS_UNCONNECTED__611, 
        SYNOPSYS_UNCONNECTED__612, SYNOPSYS_UNCONNECTED__613, \mux_out[3][31] , 
        \mux_out[3][30] , \mux_out[3][29] , \mux_out[3][28] , \mux_out[3][27] , 
        \mux_out[3][26] , \mux_out[3][25] , \mux_out[3][24] , \mux_out[3][23] , 
        \mux_out[3][22] , \mux_out[3][21] , \mux_out[3][20] , \mux_out[3][19] , 
        \mux_out[3][18] , \mux_out[3][17] , \mux_out[3][16] , \mux_out[3][15] , 
        \mux_out[3][14] , \mux_out[3][13] , \mux_out[3][12] , \mux_out[3][11] , 
        \mux_out[3][10] , \mux_out[3][9] , \mux_out[3][8] , \mux_out[3][7] , 
        \mux_out[3][6] , SYNOPSYS_UNCONNECTED__614, SYNOPSYS_UNCONNECTED__615, 
        SYNOPSYS_UNCONNECTED__616, SYNOPSYS_UNCONNECTED__617, 
        SYNOPSYS_UNCONNECTED__618, SYNOPSYS_UNCONNECTED__619}) );
  MUX_8to1_N64_12 mux_4 ( .IN0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \sub_x_1/B[23] , \sub_x_1/B[22] , 
        \sub_x_1/B[21] , A[20:18], \sub_x_1/B[17] , A[16], \sub_x_1/B[15] , 
        A[14:12], n643, n642, A[9], n641, n640, n639, n638, n637, n626, n625, 
        n636, n635, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN2({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n57, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .IN3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN4({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n32, n53, n33, n95, 
        n41, n93, n90, n50, n52, n92, n55, n96, n94, n54, n633, n631, n17, 
        n629, n19, n23, n18, n628, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .IN5({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN6({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .IN7({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .SEL({
        \encoder_out[4][2] , \encoder_out[4][1] , \encoder_out[4][0] }), .Y({
        SYNOPSYS_UNCONNECTED__620, SYNOPSYS_UNCONNECTED__621, 
        SYNOPSYS_UNCONNECTED__622, SYNOPSYS_UNCONNECTED__623, 
        SYNOPSYS_UNCONNECTED__624, SYNOPSYS_UNCONNECTED__625, 
        SYNOPSYS_UNCONNECTED__626, SYNOPSYS_UNCONNECTED__627, 
        SYNOPSYS_UNCONNECTED__628, SYNOPSYS_UNCONNECTED__629, 
        SYNOPSYS_UNCONNECTED__630, SYNOPSYS_UNCONNECTED__631, 
        SYNOPSYS_UNCONNECTED__632, SYNOPSYS_UNCONNECTED__633, 
        SYNOPSYS_UNCONNECTED__634, SYNOPSYS_UNCONNECTED__635, 
        SYNOPSYS_UNCONNECTED__636, SYNOPSYS_UNCONNECTED__637, 
        SYNOPSYS_UNCONNECTED__638, SYNOPSYS_UNCONNECTED__639, 
        SYNOPSYS_UNCONNECTED__640, SYNOPSYS_UNCONNECTED__641, 
        SYNOPSYS_UNCONNECTED__642, SYNOPSYS_UNCONNECTED__643, 
        SYNOPSYS_UNCONNECTED__644, SYNOPSYS_UNCONNECTED__645, 
        SYNOPSYS_UNCONNECTED__646, SYNOPSYS_UNCONNECTED__647, 
        SYNOPSYS_UNCONNECTED__648, SYNOPSYS_UNCONNECTED__649, 
        SYNOPSYS_UNCONNECTED__650, SYNOPSYS_UNCONNECTED__651, \mux_out[4][31] , 
        \mux_out[4][30] , \mux_out[4][29] , \mux_out[4][28] , \mux_out[4][27] , 
        \mux_out[4][26] , \mux_out[4][25] , \mux_out[4][24] , \mux_out[4][23] , 
        \mux_out[4][22] , \mux_out[4][21] , \mux_out[4][20] , \mux_out[4][19] , 
        \mux_out[4][18] , \mux_out[4][17] , \mux_out[4][16] , \mux_out[4][15] , 
        \mux_out[4][14] , \mux_out[4][13] , \mux_out[4][12] , \mux_out[4][11] , 
        \mux_out[4][10] , \mux_out[4][9] , \mux_out[4][8] , 
        SYNOPSYS_UNCONNECTED__652, SYNOPSYS_UNCONNECTED__653, 
        SYNOPSYS_UNCONNECTED__654, SYNOPSYS_UNCONNECTED__655, 
        SYNOPSYS_UNCONNECTED__656, SYNOPSYS_UNCONNECTED__657, 
        SYNOPSYS_UNCONNECTED__658, SYNOPSYS_UNCONNECTED__659}) );
  MUX_8to1_N64_11 mux_5 ( .IN0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \sub_x_1/B[21] , A[20:18], 
        \sub_x_1/B[17] , A[16], \sub_x_1/B[15] , A[14:12], n643, n642, A[9], 
        n641, n640, n639, n638, n637, n626, n625, n636, n635, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n53, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .IN3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN4({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n33, n95, n41, n93, n90, n50, n52, n91, 
        \A_shifted[-32][43] , \A_shifted[-32][42] , \A_shifted[-32][41] , 
        \A_shifted[-32][40] , n633, n632, n17, n630, n19, n23, n18, n628, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .IN5({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN6({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .IN7({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .SEL({\encoder_out[5][2] , 
        \encoder_out[5][1] , \encoder_out[5][0] }), .Y({
        SYNOPSYS_UNCONNECTED__660, SYNOPSYS_UNCONNECTED__661, 
        SYNOPSYS_UNCONNECTED__662, SYNOPSYS_UNCONNECTED__663, 
        SYNOPSYS_UNCONNECTED__664, SYNOPSYS_UNCONNECTED__665, 
        SYNOPSYS_UNCONNECTED__666, SYNOPSYS_UNCONNECTED__667, 
        SYNOPSYS_UNCONNECTED__668, SYNOPSYS_UNCONNECTED__669, 
        SYNOPSYS_UNCONNECTED__670, SYNOPSYS_UNCONNECTED__671, 
        SYNOPSYS_UNCONNECTED__672, SYNOPSYS_UNCONNECTED__673, 
        SYNOPSYS_UNCONNECTED__674, SYNOPSYS_UNCONNECTED__675, 
        SYNOPSYS_UNCONNECTED__676, SYNOPSYS_UNCONNECTED__677, 
        SYNOPSYS_UNCONNECTED__678, SYNOPSYS_UNCONNECTED__679, 
        SYNOPSYS_UNCONNECTED__680, SYNOPSYS_UNCONNECTED__681, 
        SYNOPSYS_UNCONNECTED__682, SYNOPSYS_UNCONNECTED__683, 
        SYNOPSYS_UNCONNECTED__684, SYNOPSYS_UNCONNECTED__685, 
        SYNOPSYS_UNCONNECTED__686, SYNOPSYS_UNCONNECTED__687, 
        SYNOPSYS_UNCONNECTED__688, SYNOPSYS_UNCONNECTED__689, 
        SYNOPSYS_UNCONNECTED__690, SYNOPSYS_UNCONNECTED__691, \mux_out[5][31] , 
        \mux_out[5][30] , \mux_out[5][29] , \mux_out[5][28] , \mux_out[5][27] , 
        \mux_out[5][26] , \mux_out[5][25] , \mux_out[5][24] , \mux_out[5][23] , 
        \mux_out[5][22] , \mux_out[5][21] , n22, \mux_out[5][19] , 
        \mux_out[5][18] , \mux_out[5][17] , \mux_out[5][16] , \mux_out[5][15] , 
        \mux_out[5][14] , \mux_out[5][13] , \mux_out[5][12] , \mux_out[5][11] , 
        \mux_out[5][10] , SYNOPSYS_UNCONNECTED__692, SYNOPSYS_UNCONNECTED__693, 
        SYNOPSYS_UNCONNECTED__694, SYNOPSYS_UNCONNECTED__695, 
        SYNOPSYS_UNCONNECTED__696, SYNOPSYS_UNCONNECTED__697, 
        SYNOPSYS_UNCONNECTED__698, SYNOPSYS_UNCONNECTED__699, 
        SYNOPSYS_UNCONNECTED__700, SYNOPSYS_UNCONNECTED__701}) );
  MUX_8to1_N64_10 mux_6 ( .IN0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, A[19:18], \sub_x_1/B[17] , A[16], 
        \sub_x_1/B[15] , A[14:12], n643, n642, A[9], n641, n640, n639, n638, 
        n637, n627, n625, n636, n635, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, n95, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .IN3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN4({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, n41, n93, n90, n50, n52, n92, n55, n96, n94, n54, 
        n633, n632, n17, n630, n19, n23, n18, n628, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN5({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .IN6({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN7({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .SEL({\encoder_out[6][2] , 
        \encoder_out[6][1] , \encoder_out[6][0] }), .Y({
        SYNOPSYS_UNCONNECTED__702, SYNOPSYS_UNCONNECTED__703, 
        SYNOPSYS_UNCONNECTED__704, SYNOPSYS_UNCONNECTED__705, 
        SYNOPSYS_UNCONNECTED__706, SYNOPSYS_UNCONNECTED__707, 
        SYNOPSYS_UNCONNECTED__708, SYNOPSYS_UNCONNECTED__709, 
        SYNOPSYS_UNCONNECTED__710, SYNOPSYS_UNCONNECTED__711, 
        SYNOPSYS_UNCONNECTED__712, SYNOPSYS_UNCONNECTED__713, 
        SYNOPSYS_UNCONNECTED__714, SYNOPSYS_UNCONNECTED__715, 
        SYNOPSYS_UNCONNECTED__716, SYNOPSYS_UNCONNECTED__717, 
        SYNOPSYS_UNCONNECTED__718, SYNOPSYS_UNCONNECTED__719, 
        SYNOPSYS_UNCONNECTED__720, SYNOPSYS_UNCONNECTED__721, 
        SYNOPSYS_UNCONNECTED__722, SYNOPSYS_UNCONNECTED__723, 
        SYNOPSYS_UNCONNECTED__724, SYNOPSYS_UNCONNECTED__725, 
        SYNOPSYS_UNCONNECTED__726, SYNOPSYS_UNCONNECTED__727, 
        SYNOPSYS_UNCONNECTED__728, SYNOPSYS_UNCONNECTED__729, 
        SYNOPSYS_UNCONNECTED__730, SYNOPSYS_UNCONNECTED__731, 
        SYNOPSYS_UNCONNECTED__732, SYNOPSYS_UNCONNECTED__733, \mux_out[6][31] , 
        \mux_out[6][30] , \mux_out[6][29] , \mux_out[6][28] , \mux_out[6][27] , 
        \mux_out[6][26] , \mux_out[6][25] , \mux_out[6][24] , \mux_out[6][23] , 
        \mux_out[6][22] , \mux_out[6][21] , \mux_out[6][20] , \mux_out[6][19] , 
        \mux_out[6][18] , \mux_out[6][17] , \mux_out[6][16] , \mux_out[6][15] , 
        \mux_out[6][14] , \mux_out[6][13] , \mux_out[6][12] , 
        SYNOPSYS_UNCONNECTED__734, SYNOPSYS_UNCONNECTED__735, 
        SYNOPSYS_UNCONNECTED__736, SYNOPSYS_UNCONNECTED__737, 
        SYNOPSYS_UNCONNECTED__738, SYNOPSYS_UNCONNECTED__739, 
        SYNOPSYS_UNCONNECTED__740, SYNOPSYS_UNCONNECTED__741, 
        SYNOPSYS_UNCONNECTED__742, SYNOPSYS_UNCONNECTED__743, 
        SYNOPSYS_UNCONNECTED__744, SYNOPSYS_UNCONNECTED__745}) );
  MUX_8to1_N64_9 mux_7 ( .IN0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \sub_x_1/B[17] , A[16], 
        \sub_x_1/B[15] , A[14:12], n643, n642, A[9], n641, n640, n639, n638, 
        n637, n626, n625, n636, n635, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN2({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n93, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .IN3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN4({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n90, n50, n52, n92, n55, n96, n94, n54, 
        n633, n631, n17, n629, n19, n23, n18, n628, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN5({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN6({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .IN7({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .SEL({\encoder_out[7][2] , 
        \encoder_out[7][1] , \encoder_out[7][0] }), .Y({
        SYNOPSYS_UNCONNECTED__746, SYNOPSYS_UNCONNECTED__747, 
        SYNOPSYS_UNCONNECTED__748, SYNOPSYS_UNCONNECTED__749, 
        SYNOPSYS_UNCONNECTED__750, SYNOPSYS_UNCONNECTED__751, 
        SYNOPSYS_UNCONNECTED__752, SYNOPSYS_UNCONNECTED__753, 
        SYNOPSYS_UNCONNECTED__754, SYNOPSYS_UNCONNECTED__755, 
        SYNOPSYS_UNCONNECTED__756, SYNOPSYS_UNCONNECTED__757, 
        SYNOPSYS_UNCONNECTED__758, SYNOPSYS_UNCONNECTED__759, 
        SYNOPSYS_UNCONNECTED__760, SYNOPSYS_UNCONNECTED__761, 
        SYNOPSYS_UNCONNECTED__762, SYNOPSYS_UNCONNECTED__763, 
        SYNOPSYS_UNCONNECTED__764, SYNOPSYS_UNCONNECTED__765, 
        SYNOPSYS_UNCONNECTED__766, SYNOPSYS_UNCONNECTED__767, 
        SYNOPSYS_UNCONNECTED__768, SYNOPSYS_UNCONNECTED__769, 
        SYNOPSYS_UNCONNECTED__770, SYNOPSYS_UNCONNECTED__771, 
        SYNOPSYS_UNCONNECTED__772, SYNOPSYS_UNCONNECTED__773, 
        SYNOPSYS_UNCONNECTED__774, SYNOPSYS_UNCONNECTED__775, 
        SYNOPSYS_UNCONNECTED__776, SYNOPSYS_UNCONNECTED__777, \mux_out[7][31] , 
        \mux_out[7][30] , \mux_out[7][29] , \mux_out[7][28] , \mux_out[7][27] , 
        \mux_out[7][26] , \mux_out[7][25] , \mux_out[7][24] , \mux_out[7][23] , 
        \mux_out[7][22] , \mux_out[7][21] , \mux_out[7][20] , \mux_out[7][19] , 
        \mux_out[7][18] , \mux_out[7][17] , \mux_out[7][16] , \mux_out[7][15] , 
        \mux_out[7][14] , SYNOPSYS_UNCONNECTED__778, SYNOPSYS_UNCONNECTED__779, 
        SYNOPSYS_UNCONNECTED__780, SYNOPSYS_UNCONNECTED__781, 
        SYNOPSYS_UNCONNECTED__782, SYNOPSYS_UNCONNECTED__783, 
        SYNOPSYS_UNCONNECTED__784, SYNOPSYS_UNCONNECTED__785, 
        SYNOPSYS_UNCONNECTED__786, SYNOPSYS_UNCONNECTED__787, 
        SYNOPSYS_UNCONNECTED__788, SYNOPSYS_UNCONNECTED__789, 
        SYNOPSYS_UNCONNECTED__790, SYNOPSYS_UNCONNECTED__791}) );
  MUX_8to1_N64_8 mux_8 ( .IN0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \sub_x_1/B[15] , A[14:12], n643, 
        n642, A[9], n641, n640, n639, A[5], n637, n626, n625, n636, n635, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .IN2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, n50, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN3({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .IN4({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, n52, n92, n55, n96, n94, n54, n634, n631, n17, n629, n19, n23, 
        n18, n628, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN5({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .IN6({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN7({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .SEL({\encoder_out[8][2] , \encoder_out[8][1] , 
        \encoder_out[8][0] }), .Y({SYNOPSYS_UNCONNECTED__792, 
        SYNOPSYS_UNCONNECTED__793, SYNOPSYS_UNCONNECTED__794, 
        SYNOPSYS_UNCONNECTED__795, SYNOPSYS_UNCONNECTED__796, 
        SYNOPSYS_UNCONNECTED__797, SYNOPSYS_UNCONNECTED__798, 
        SYNOPSYS_UNCONNECTED__799, SYNOPSYS_UNCONNECTED__800, 
        SYNOPSYS_UNCONNECTED__801, SYNOPSYS_UNCONNECTED__802, 
        SYNOPSYS_UNCONNECTED__803, SYNOPSYS_UNCONNECTED__804, 
        SYNOPSYS_UNCONNECTED__805, SYNOPSYS_UNCONNECTED__806, 
        SYNOPSYS_UNCONNECTED__807, SYNOPSYS_UNCONNECTED__808, 
        SYNOPSYS_UNCONNECTED__809, SYNOPSYS_UNCONNECTED__810, 
        SYNOPSYS_UNCONNECTED__811, SYNOPSYS_UNCONNECTED__812, 
        SYNOPSYS_UNCONNECTED__813, SYNOPSYS_UNCONNECTED__814, 
        SYNOPSYS_UNCONNECTED__815, SYNOPSYS_UNCONNECTED__816, 
        SYNOPSYS_UNCONNECTED__817, SYNOPSYS_UNCONNECTED__818, 
        SYNOPSYS_UNCONNECTED__819, SYNOPSYS_UNCONNECTED__820, 
        SYNOPSYS_UNCONNECTED__821, SYNOPSYS_UNCONNECTED__822, 
        SYNOPSYS_UNCONNECTED__823, \mux_out[8][31] , \mux_out[8][30] , 
        \mux_out[8][29] , \mux_out[8][28] , \mux_out[8][27] , \mux_out[8][26] , 
        \mux_out[8][25] , \mux_out[8][24] , \mux_out[8][23] , \mux_out[8][22] , 
        \mux_out[8][21] , \mux_out[8][20] , \mux_out[8][19] , \mux_out[8][18] , 
        \mux_out[8][17] , \mux_out[8][16] , SYNOPSYS_UNCONNECTED__824, 
        SYNOPSYS_UNCONNECTED__825, SYNOPSYS_UNCONNECTED__826, 
        SYNOPSYS_UNCONNECTED__827, SYNOPSYS_UNCONNECTED__828, 
        SYNOPSYS_UNCONNECTED__829, SYNOPSYS_UNCONNECTED__830, 
        SYNOPSYS_UNCONNECTED__831, SYNOPSYS_UNCONNECTED__832, 
        SYNOPSYS_UNCONNECTED__833, SYNOPSYS_UNCONNECTED__834, 
        SYNOPSYS_UNCONNECTED__835, SYNOPSYS_UNCONNECTED__836, 
        SYNOPSYS_UNCONNECTED__837, SYNOPSYS_UNCONNECTED__838, 
        SYNOPSYS_UNCONNECTED__839}) );
  MUX_8to1_N64_7 mux_9 ( .IN0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, A[13:12], n643, n642, A[9], n641, 
        n640, n639, n638, n637, n626, n625, n636, n635, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .IN2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        n92, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN3({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .IN4({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        n55, n96, n94, n54, n633, n631, n17, n629, n19, n23, n18, n628, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN5({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .IN6({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN7({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .SEL({\encoder_out[9][2] , \encoder_out[9][1] , 
        \encoder_out[9][0] }), .Y({SYNOPSYS_UNCONNECTED__840, 
        SYNOPSYS_UNCONNECTED__841, SYNOPSYS_UNCONNECTED__842, 
        SYNOPSYS_UNCONNECTED__843, SYNOPSYS_UNCONNECTED__844, 
        SYNOPSYS_UNCONNECTED__845, SYNOPSYS_UNCONNECTED__846, 
        SYNOPSYS_UNCONNECTED__847, SYNOPSYS_UNCONNECTED__848, 
        SYNOPSYS_UNCONNECTED__849, SYNOPSYS_UNCONNECTED__850, 
        SYNOPSYS_UNCONNECTED__851, SYNOPSYS_UNCONNECTED__852, 
        SYNOPSYS_UNCONNECTED__853, SYNOPSYS_UNCONNECTED__854, 
        SYNOPSYS_UNCONNECTED__855, SYNOPSYS_UNCONNECTED__856, 
        SYNOPSYS_UNCONNECTED__857, SYNOPSYS_UNCONNECTED__858, 
        SYNOPSYS_UNCONNECTED__859, SYNOPSYS_UNCONNECTED__860, 
        SYNOPSYS_UNCONNECTED__861, SYNOPSYS_UNCONNECTED__862, 
        SYNOPSYS_UNCONNECTED__863, SYNOPSYS_UNCONNECTED__864, 
        SYNOPSYS_UNCONNECTED__865, SYNOPSYS_UNCONNECTED__866, 
        SYNOPSYS_UNCONNECTED__867, SYNOPSYS_UNCONNECTED__868, 
        SYNOPSYS_UNCONNECTED__869, SYNOPSYS_UNCONNECTED__870, 
        SYNOPSYS_UNCONNECTED__871, \mux_out[9][31] , \mux_out[9][30] , 
        \mux_out[9][29] , \mux_out[9][28] , \mux_out[9][27] , \mux_out[9][26] , 
        \mux_out[9][25] , \mux_out[9][24] , \mux_out[9][23] , \mux_out[9][22] , 
        \mux_out[9][21] , \mux_out[9][20] , \mux_out[9][19] , \mux_out[9][18] , 
        SYNOPSYS_UNCONNECTED__872, SYNOPSYS_UNCONNECTED__873, 
        SYNOPSYS_UNCONNECTED__874, SYNOPSYS_UNCONNECTED__875, 
        SYNOPSYS_UNCONNECTED__876, SYNOPSYS_UNCONNECTED__877, 
        SYNOPSYS_UNCONNECTED__878, SYNOPSYS_UNCONNECTED__879, 
        SYNOPSYS_UNCONNECTED__880, SYNOPSYS_UNCONNECTED__881, 
        SYNOPSYS_UNCONNECTED__882, SYNOPSYS_UNCONNECTED__883, 
        SYNOPSYS_UNCONNECTED__884, SYNOPSYS_UNCONNECTED__885, 
        SYNOPSYS_UNCONNECTED__886, SYNOPSYS_UNCONNECTED__887, 
        SYNOPSYS_UNCONNECTED__888, SYNOPSYS_UNCONNECTED__889}) );
  MUX_8to1_N64_6 mux_10 ( .IN0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n643, n642, A[9], n641, n640, n639, 
        n638, n637, n627, n625, n636, n635, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .IN2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        n96, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN3({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .IN4({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        n94, n54, n634, n631, n17, n629, n19, n23, n18, n628, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN5({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .IN6({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN7({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .SEL({\encoder_out[10][2] , \encoder_out[10][1] , 
        \encoder_out[10][0] }), .Y({SYNOPSYS_UNCONNECTED__890, 
        SYNOPSYS_UNCONNECTED__891, SYNOPSYS_UNCONNECTED__892, 
        SYNOPSYS_UNCONNECTED__893, SYNOPSYS_UNCONNECTED__894, 
        SYNOPSYS_UNCONNECTED__895, SYNOPSYS_UNCONNECTED__896, 
        SYNOPSYS_UNCONNECTED__897, SYNOPSYS_UNCONNECTED__898, 
        SYNOPSYS_UNCONNECTED__899, SYNOPSYS_UNCONNECTED__900, 
        SYNOPSYS_UNCONNECTED__901, SYNOPSYS_UNCONNECTED__902, 
        SYNOPSYS_UNCONNECTED__903, SYNOPSYS_UNCONNECTED__904, 
        SYNOPSYS_UNCONNECTED__905, SYNOPSYS_UNCONNECTED__906, 
        SYNOPSYS_UNCONNECTED__907, SYNOPSYS_UNCONNECTED__908, 
        SYNOPSYS_UNCONNECTED__909, SYNOPSYS_UNCONNECTED__910, 
        SYNOPSYS_UNCONNECTED__911, SYNOPSYS_UNCONNECTED__912, 
        SYNOPSYS_UNCONNECTED__913, SYNOPSYS_UNCONNECTED__914, 
        SYNOPSYS_UNCONNECTED__915, SYNOPSYS_UNCONNECTED__916, 
        SYNOPSYS_UNCONNECTED__917, SYNOPSYS_UNCONNECTED__918, 
        SYNOPSYS_UNCONNECTED__919, SYNOPSYS_UNCONNECTED__920, 
        SYNOPSYS_UNCONNECTED__921, \mux_out[10][31] , \mux_out[10][30] , 
        \mux_out[10][29] , \mux_out[10][28] , \mux_out[10][27] , 
        \mux_out[10][26] , \mux_out[10][25] , \mux_out[10][24] , 
        \mux_out[10][23] , \mux_out[10][22] , \mux_out[10][21] , 
        \mux_out[10][20] , SYNOPSYS_UNCONNECTED__922, 
        SYNOPSYS_UNCONNECTED__923, SYNOPSYS_UNCONNECTED__924, 
        SYNOPSYS_UNCONNECTED__925, SYNOPSYS_UNCONNECTED__926, 
        SYNOPSYS_UNCONNECTED__927, SYNOPSYS_UNCONNECTED__928, 
        SYNOPSYS_UNCONNECTED__929, SYNOPSYS_UNCONNECTED__930, 
        SYNOPSYS_UNCONNECTED__931, SYNOPSYS_UNCONNECTED__932, 
        SYNOPSYS_UNCONNECTED__933, SYNOPSYS_UNCONNECTED__934, 
        SYNOPSYS_UNCONNECTED__935, SYNOPSYS_UNCONNECTED__936, 
        SYNOPSYS_UNCONNECTED__937, SYNOPSYS_UNCONNECTED__938, 
        SYNOPSYS_UNCONNECTED__939, SYNOPSYS_UNCONNECTED__940, 
        SYNOPSYS_UNCONNECTED__941}) );
  MUX_8to1_N64_5 mux_11 ( .IN0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, A[9], n641, n640, n639, n638, n637, 
        n627, n625, n636, n635, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .IN2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        n54, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN3({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .IN4({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        n633, n631, n17, n629, n19, n23, n18, n628, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN5({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .IN6({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN7({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .SEL({\encoder_out[11][2] , \encoder_out[11][1] , 
        \encoder_out[11][0] }), .Y({SYNOPSYS_UNCONNECTED__942, 
        SYNOPSYS_UNCONNECTED__943, SYNOPSYS_UNCONNECTED__944, 
        SYNOPSYS_UNCONNECTED__945, SYNOPSYS_UNCONNECTED__946, 
        SYNOPSYS_UNCONNECTED__947, SYNOPSYS_UNCONNECTED__948, 
        SYNOPSYS_UNCONNECTED__949, SYNOPSYS_UNCONNECTED__950, 
        SYNOPSYS_UNCONNECTED__951, SYNOPSYS_UNCONNECTED__952, 
        SYNOPSYS_UNCONNECTED__953, SYNOPSYS_UNCONNECTED__954, 
        SYNOPSYS_UNCONNECTED__955, SYNOPSYS_UNCONNECTED__956, 
        SYNOPSYS_UNCONNECTED__957, SYNOPSYS_UNCONNECTED__958, 
        SYNOPSYS_UNCONNECTED__959, SYNOPSYS_UNCONNECTED__960, 
        SYNOPSYS_UNCONNECTED__961, SYNOPSYS_UNCONNECTED__962, 
        SYNOPSYS_UNCONNECTED__963, SYNOPSYS_UNCONNECTED__964, 
        SYNOPSYS_UNCONNECTED__965, SYNOPSYS_UNCONNECTED__966, 
        SYNOPSYS_UNCONNECTED__967, SYNOPSYS_UNCONNECTED__968, 
        SYNOPSYS_UNCONNECTED__969, SYNOPSYS_UNCONNECTED__970, 
        SYNOPSYS_UNCONNECTED__971, SYNOPSYS_UNCONNECTED__972, 
        SYNOPSYS_UNCONNECTED__973, \mux_out[11][31] , \mux_out[11][30] , 
        \mux_out[11][29] , \mux_out[11][28] , \mux_out[11][27] , 
        \mux_out[11][26] , \mux_out[11][25] , \mux_out[11][24] , 
        \mux_out[11][23] , \mux_out[11][22] , SYNOPSYS_UNCONNECTED__974, 
        SYNOPSYS_UNCONNECTED__975, SYNOPSYS_UNCONNECTED__976, 
        SYNOPSYS_UNCONNECTED__977, SYNOPSYS_UNCONNECTED__978, 
        SYNOPSYS_UNCONNECTED__979, SYNOPSYS_UNCONNECTED__980, 
        SYNOPSYS_UNCONNECTED__981, SYNOPSYS_UNCONNECTED__982, 
        SYNOPSYS_UNCONNECTED__983, SYNOPSYS_UNCONNECTED__984, 
        SYNOPSYS_UNCONNECTED__985, SYNOPSYS_UNCONNECTED__986, 
        SYNOPSYS_UNCONNECTED__987, SYNOPSYS_UNCONNECTED__988, 
        SYNOPSYS_UNCONNECTED__989, SYNOPSYS_UNCONNECTED__990, 
        SYNOPSYS_UNCONNECTED__991, SYNOPSYS_UNCONNECTED__992, 
        SYNOPSYS_UNCONNECTED__993, SYNOPSYS_UNCONNECTED__994, 
        SYNOPSYS_UNCONNECTED__995}) );
  MUX_8to1_N64_4 mux_12 ( .IN0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n640, A[6], n638, n637, n627, n625, 
        n636, n635, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .IN2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        n632, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN3({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .IN4({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        n17, n629, n19, n23, n18, n628, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN5({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .IN6({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN7({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .SEL({\encoder_out[12][2] , \encoder_out[12][1] , 
        \encoder_out[12][0] }), .Y({SYNOPSYS_UNCONNECTED__996, 
        SYNOPSYS_UNCONNECTED__997, SYNOPSYS_UNCONNECTED__998, 
        SYNOPSYS_UNCONNECTED__999, SYNOPSYS_UNCONNECTED__1000, 
        SYNOPSYS_UNCONNECTED__1001, SYNOPSYS_UNCONNECTED__1002, 
        SYNOPSYS_UNCONNECTED__1003, SYNOPSYS_UNCONNECTED__1004, 
        SYNOPSYS_UNCONNECTED__1005, SYNOPSYS_UNCONNECTED__1006, 
        SYNOPSYS_UNCONNECTED__1007, SYNOPSYS_UNCONNECTED__1008, 
        SYNOPSYS_UNCONNECTED__1009, SYNOPSYS_UNCONNECTED__1010, 
        SYNOPSYS_UNCONNECTED__1011, SYNOPSYS_UNCONNECTED__1012, 
        SYNOPSYS_UNCONNECTED__1013, SYNOPSYS_UNCONNECTED__1014, 
        SYNOPSYS_UNCONNECTED__1015, SYNOPSYS_UNCONNECTED__1016, 
        SYNOPSYS_UNCONNECTED__1017, SYNOPSYS_UNCONNECTED__1018, 
        SYNOPSYS_UNCONNECTED__1019, SYNOPSYS_UNCONNECTED__1020, 
        SYNOPSYS_UNCONNECTED__1021, SYNOPSYS_UNCONNECTED__1022, 
        SYNOPSYS_UNCONNECTED__1023, SYNOPSYS_UNCONNECTED__1024, 
        SYNOPSYS_UNCONNECTED__1025, SYNOPSYS_UNCONNECTED__1026, 
        SYNOPSYS_UNCONNECTED__1027, \mux_out[12][31] , \mux_out[12][30] , 
        \mux_out[12][29] , \mux_out[12][28] , \mux_out[12][27] , 
        \mux_out[12][26] , \mux_out[12][25] , \mux_out[12][24] , 
        SYNOPSYS_UNCONNECTED__1028, SYNOPSYS_UNCONNECTED__1029, 
        SYNOPSYS_UNCONNECTED__1030, SYNOPSYS_UNCONNECTED__1031, 
        SYNOPSYS_UNCONNECTED__1032, SYNOPSYS_UNCONNECTED__1033, 
        SYNOPSYS_UNCONNECTED__1034, SYNOPSYS_UNCONNECTED__1035, 
        SYNOPSYS_UNCONNECTED__1036, SYNOPSYS_UNCONNECTED__1037, 
        SYNOPSYS_UNCONNECTED__1038, SYNOPSYS_UNCONNECTED__1039, 
        SYNOPSYS_UNCONNECTED__1040, SYNOPSYS_UNCONNECTED__1041, 
        SYNOPSYS_UNCONNECTED__1042, SYNOPSYS_UNCONNECTED__1043, 
        SYNOPSYS_UNCONNECTED__1044, SYNOPSYS_UNCONNECTED__1045, 
        SYNOPSYS_UNCONNECTED__1046, SYNOPSYS_UNCONNECTED__1047, 
        SYNOPSYS_UNCONNECTED__1048, SYNOPSYS_UNCONNECTED__1049, 
        SYNOPSYS_UNCONNECTED__1050, SYNOPSYS_UNCONNECTED__1051}) );
  MUX_8to1_N64_3 mux_13 ( .IN0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n638, n637, n627, n625, n636, n635, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .IN2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        n630, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN3({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .IN4({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        n19, n23, n18, n628, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN5({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .IN6({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN7({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .SEL({\encoder_out[13][2] , \encoder_out[13][1] , 
        \encoder_out[13][0] }), .Y({SYNOPSYS_UNCONNECTED__1052, 
        SYNOPSYS_UNCONNECTED__1053, SYNOPSYS_UNCONNECTED__1054, 
        SYNOPSYS_UNCONNECTED__1055, SYNOPSYS_UNCONNECTED__1056, 
        SYNOPSYS_UNCONNECTED__1057, SYNOPSYS_UNCONNECTED__1058, 
        SYNOPSYS_UNCONNECTED__1059, SYNOPSYS_UNCONNECTED__1060, 
        SYNOPSYS_UNCONNECTED__1061, SYNOPSYS_UNCONNECTED__1062, 
        SYNOPSYS_UNCONNECTED__1063, SYNOPSYS_UNCONNECTED__1064, 
        SYNOPSYS_UNCONNECTED__1065, SYNOPSYS_UNCONNECTED__1066, 
        SYNOPSYS_UNCONNECTED__1067, SYNOPSYS_UNCONNECTED__1068, 
        SYNOPSYS_UNCONNECTED__1069, SYNOPSYS_UNCONNECTED__1070, 
        SYNOPSYS_UNCONNECTED__1071, SYNOPSYS_UNCONNECTED__1072, 
        SYNOPSYS_UNCONNECTED__1073, SYNOPSYS_UNCONNECTED__1074, 
        SYNOPSYS_UNCONNECTED__1075, SYNOPSYS_UNCONNECTED__1076, 
        SYNOPSYS_UNCONNECTED__1077, SYNOPSYS_UNCONNECTED__1078, 
        SYNOPSYS_UNCONNECTED__1079, SYNOPSYS_UNCONNECTED__1080, 
        SYNOPSYS_UNCONNECTED__1081, SYNOPSYS_UNCONNECTED__1082, 
        SYNOPSYS_UNCONNECTED__1083, \mux_out[13][31] , \mux_out[13][30] , 
        \mux_out[13][29] , \mux_out[13][28] , \mux_out[13][27] , 
        \mux_out[13][26] , SYNOPSYS_UNCONNECTED__1084, 
        SYNOPSYS_UNCONNECTED__1085, SYNOPSYS_UNCONNECTED__1086, 
        SYNOPSYS_UNCONNECTED__1087, SYNOPSYS_UNCONNECTED__1088, 
        SYNOPSYS_UNCONNECTED__1089, SYNOPSYS_UNCONNECTED__1090, 
        SYNOPSYS_UNCONNECTED__1091, SYNOPSYS_UNCONNECTED__1092, 
        SYNOPSYS_UNCONNECTED__1093, SYNOPSYS_UNCONNECTED__1094, 
        SYNOPSYS_UNCONNECTED__1095, SYNOPSYS_UNCONNECTED__1096, 
        SYNOPSYS_UNCONNECTED__1097, SYNOPSYS_UNCONNECTED__1098, 
        SYNOPSYS_UNCONNECTED__1099, SYNOPSYS_UNCONNECTED__1100, 
        SYNOPSYS_UNCONNECTED__1101, SYNOPSYS_UNCONNECTED__1102, 
        SYNOPSYS_UNCONNECTED__1103, SYNOPSYS_UNCONNECTED__1104, 
        SYNOPSYS_UNCONNECTED__1105, SYNOPSYS_UNCONNECTED__1106, 
        SYNOPSYS_UNCONNECTED__1107, SYNOPSYS_UNCONNECTED__1108, 
        SYNOPSYS_UNCONNECTED__1109}) );
  MUX_8to1_N64_2 mux_14 ( .IN0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n627, n625, n636, n635, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .IN2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        n23, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN3({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .IN4({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        n18, n628, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN5({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .IN6({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN7({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .SEL({\encoder_out[14][2] , \encoder_out[14][1] , 
        \encoder_out[14][0] }), .Y({SYNOPSYS_UNCONNECTED__1110, 
        SYNOPSYS_UNCONNECTED__1111, SYNOPSYS_UNCONNECTED__1112, 
        SYNOPSYS_UNCONNECTED__1113, SYNOPSYS_UNCONNECTED__1114, 
        SYNOPSYS_UNCONNECTED__1115, SYNOPSYS_UNCONNECTED__1116, 
        SYNOPSYS_UNCONNECTED__1117, SYNOPSYS_UNCONNECTED__1118, 
        SYNOPSYS_UNCONNECTED__1119, SYNOPSYS_UNCONNECTED__1120, 
        SYNOPSYS_UNCONNECTED__1121, SYNOPSYS_UNCONNECTED__1122, 
        SYNOPSYS_UNCONNECTED__1123, SYNOPSYS_UNCONNECTED__1124, 
        SYNOPSYS_UNCONNECTED__1125, SYNOPSYS_UNCONNECTED__1126, 
        SYNOPSYS_UNCONNECTED__1127, SYNOPSYS_UNCONNECTED__1128, 
        SYNOPSYS_UNCONNECTED__1129, SYNOPSYS_UNCONNECTED__1130, 
        SYNOPSYS_UNCONNECTED__1131, SYNOPSYS_UNCONNECTED__1132, 
        SYNOPSYS_UNCONNECTED__1133, SYNOPSYS_UNCONNECTED__1134, 
        SYNOPSYS_UNCONNECTED__1135, SYNOPSYS_UNCONNECTED__1136, 
        SYNOPSYS_UNCONNECTED__1137, SYNOPSYS_UNCONNECTED__1138, 
        SYNOPSYS_UNCONNECTED__1139, SYNOPSYS_UNCONNECTED__1140, 
        SYNOPSYS_UNCONNECTED__1141, \mux_out[14][31] , \mux_out[14][30] , 
        \mux_out[14][29] , \mux_out[14][28] , SYNOPSYS_UNCONNECTED__1142, 
        SYNOPSYS_UNCONNECTED__1143, SYNOPSYS_UNCONNECTED__1144, 
        SYNOPSYS_UNCONNECTED__1145, SYNOPSYS_UNCONNECTED__1146, 
        SYNOPSYS_UNCONNECTED__1147, SYNOPSYS_UNCONNECTED__1148, 
        SYNOPSYS_UNCONNECTED__1149, SYNOPSYS_UNCONNECTED__1150, 
        SYNOPSYS_UNCONNECTED__1151, SYNOPSYS_UNCONNECTED__1152, 
        SYNOPSYS_UNCONNECTED__1153, SYNOPSYS_UNCONNECTED__1154, 
        SYNOPSYS_UNCONNECTED__1155, SYNOPSYS_UNCONNECTED__1156, 
        SYNOPSYS_UNCONNECTED__1157, SYNOPSYS_UNCONNECTED__1158, 
        SYNOPSYS_UNCONNECTED__1159, SYNOPSYS_UNCONNECTED__1160, 
        SYNOPSYS_UNCONNECTED__1161, SYNOPSYS_UNCONNECTED__1162, 
        SYNOPSYS_UNCONNECTED__1163, SYNOPSYS_UNCONNECTED__1164, 
        SYNOPSYS_UNCONNECTED__1165, SYNOPSYS_UNCONNECTED__1166, 
        SYNOPSYS_UNCONNECTED__1167, SYNOPSYS_UNCONNECTED__1168, 
        SYNOPSYS_UNCONNECTED__1169}) );
  MUX_8to1_N64_1 mux_15 ( .IN0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN1({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n636, n635, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .IN2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        n628, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN3({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .IN4({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN5({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .IN6({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN7({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .SEL({\encoder_out[15][2] , \encoder_out[15][1] , 
        \encoder_out[15][0] }), .Y({SYNOPSYS_UNCONNECTED__1170, 
        SYNOPSYS_UNCONNECTED__1171, SYNOPSYS_UNCONNECTED__1172, 
        SYNOPSYS_UNCONNECTED__1173, SYNOPSYS_UNCONNECTED__1174, 
        SYNOPSYS_UNCONNECTED__1175, SYNOPSYS_UNCONNECTED__1176, 
        SYNOPSYS_UNCONNECTED__1177, SYNOPSYS_UNCONNECTED__1178, 
        SYNOPSYS_UNCONNECTED__1179, SYNOPSYS_UNCONNECTED__1180, 
        SYNOPSYS_UNCONNECTED__1181, SYNOPSYS_UNCONNECTED__1182, 
        SYNOPSYS_UNCONNECTED__1183, SYNOPSYS_UNCONNECTED__1184, 
        SYNOPSYS_UNCONNECTED__1185, SYNOPSYS_UNCONNECTED__1186, 
        SYNOPSYS_UNCONNECTED__1187, SYNOPSYS_UNCONNECTED__1188, 
        SYNOPSYS_UNCONNECTED__1189, SYNOPSYS_UNCONNECTED__1190, 
        SYNOPSYS_UNCONNECTED__1191, SYNOPSYS_UNCONNECTED__1192, 
        SYNOPSYS_UNCONNECTED__1193, SYNOPSYS_UNCONNECTED__1194, 
        SYNOPSYS_UNCONNECTED__1195, SYNOPSYS_UNCONNECTED__1196, 
        SYNOPSYS_UNCONNECTED__1197, SYNOPSYS_UNCONNECTED__1198, 
        SYNOPSYS_UNCONNECTED__1199, SYNOPSYS_UNCONNECTED__1200, 
        SYNOPSYS_UNCONNECTED__1201, \mux_out[15][31] , \mux_out[15][30] , 
        SYNOPSYS_UNCONNECTED__1202, SYNOPSYS_UNCONNECTED__1203, 
        SYNOPSYS_UNCONNECTED__1204, SYNOPSYS_UNCONNECTED__1205, 
        SYNOPSYS_UNCONNECTED__1206, SYNOPSYS_UNCONNECTED__1207, 
        SYNOPSYS_UNCONNECTED__1208, SYNOPSYS_UNCONNECTED__1209, 
        SYNOPSYS_UNCONNECTED__1210, SYNOPSYS_UNCONNECTED__1211, 
        SYNOPSYS_UNCONNECTED__1212, SYNOPSYS_UNCONNECTED__1213, 
        SYNOPSYS_UNCONNECTED__1214, SYNOPSYS_UNCONNECTED__1215, 
        SYNOPSYS_UNCONNECTED__1216, SYNOPSYS_UNCONNECTED__1217, 
        SYNOPSYS_UNCONNECTED__1218, SYNOPSYS_UNCONNECTED__1219, 
        SYNOPSYS_UNCONNECTED__1220, SYNOPSYS_UNCONNECTED__1221, 
        SYNOPSYS_UNCONNECTED__1222, SYNOPSYS_UNCONNECTED__1223, 
        SYNOPSYS_UNCONNECTED__1224, SYNOPSYS_UNCONNECTED__1225, 
        SYNOPSYS_UNCONNECTED__1226, SYNOPSYS_UNCONNECTED__1227, 
        SYNOPSYS_UNCONNECTED__1228, SYNOPSYS_UNCONNECTED__1229, 
        SYNOPSYS_UNCONNECTED__1230, SYNOPSYS_UNCONNECTED__1231}) );
  booth_encoder_0 encoder_0 ( .\input ({B[1:0], 1'b0}), .\output ({
        \encoder_out[0][2] , \encoder_out[0][1] , \encoder_out[0][0] }) );
  booth_encoder_15 encoder_1 ( .\input (B[3:1]), .\output ({
        \encoder_out[1][2] , \encoder_out[1][1] , \encoder_out[1][0] }) );
  booth_encoder_14 encoder_2 ( .\input (B[5:3]), .\output ({
        \encoder_out[2][2] , \encoder_out[2][1] , \encoder_out[2][0] }) );
  booth_encoder_13 encoder_3 ( .\input (B[7:5]), .\output ({
        \encoder_out[3][2] , \encoder_out[3][1] , \encoder_out[3][0] }) );
  booth_encoder_12 encoder_4 ( .\input ({n46, B[8:7]}), .\output ({
        \encoder_out[4][2] , \encoder_out[4][1] , \encoder_out[4][0] }) );
  booth_encoder_11 encoder_5 ( .\input (B[11:9]), .\output ({
        \encoder_out[5][2] , \encoder_out[5][1] , \encoder_out[5][0] }) );
  booth_encoder_10 encoder_6 ( .\input (B[13:11]), .\output ({
        \encoder_out[6][2] , \encoder_out[6][1] , \encoder_out[6][0] }) );
  booth_encoder_9 encoder_7 ( .\input (B[15:13]), .\output ({
        \encoder_out[7][2] , \encoder_out[7][1] , \encoder_out[7][0] }) );
  booth_encoder_8 encoder_8 ( .\input (B[17:15]), .\output ({
        \encoder_out[8][2] , \encoder_out[8][1] , \encoder_out[8][0] }) );
  booth_encoder_7 encoder_9 ( .\input (B[19:17]), .\output ({
        \encoder_out[9][2] , \encoder_out[9][1] , \encoder_out[9][0] }) );
  booth_encoder_6 encoder_10 ( .\input (B[21:19]), .\output ({
        \encoder_out[10][2] , \encoder_out[10][1] , \encoder_out[10][0] }) );
  booth_encoder_5 encoder_11 ( .\input (B[23:21]), .\output ({
        \encoder_out[11][2] , \encoder_out[11][1] , \encoder_out[11][0] }) );
  booth_encoder_4 encoder_12 ( .\input ({n44, B[24:23]}), .\output ({
        \encoder_out[12][2] , \encoder_out[12][1] , \encoder_out[12][0] }) );
  booth_encoder_3 encoder_13 ( .\input (B[27:25]), .\output ({
        \encoder_out[13][2] , \encoder_out[13][1] , \encoder_out[13][0] }) );
  booth_encoder_2 encoder_14 ( .\input (B[29:27]), .\output ({
        \encoder_out[14][2] , \encoder_out[14][1] , \encoder_out[14][0] }) );
  booth_encoder_1 encoder_15 ( .\input (B[31:29]), .\output ({
        \encoder_out[15][2] , \encoder_out[15][1] , \encoder_out[15][0] }) );
  SNPS_CLOCK_GATE_HIGH_boothmul_4stage_N32_5 \clk_gate_add_out_s4_reg[12]_0  ( 
        .CLK(CLK), .EN(EN), .ENCLK(net18822), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_boothmul_4stage_N32_3 \clk_gate_add_out_s2_reg[4]_0  ( 
        .CLK(CLK), .EN(EN), .ENCLK(net18832), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_boothmul_4stage_N32_1 \clk_gate_add_out_s3_reg[8]_0  ( 
        .CLK(CLK), .EN(EN), .ENCLK(net18842), .TE(1'b0) );
  DFFR_X1 \add_out_s2_reg[4][26]  ( .D(\add_out_s1[4][26] ), .CK(net18832), 
        .RN(RST), .Q(\add_out_s2[4][26] ) );
  DFFR_X1 \add_out_s2_reg[4][25]  ( .D(\add_out_s1[4][25] ), .CK(net18832), 
        .RN(RST), .Q(\add_out_s2[4][25] ) );
  DFFR_X1 \add_out_s2_reg[4][24]  ( .D(\add_out_s1[4][24] ), .CK(net18832), 
        .RN(RST), .Q(\add_out_s2[4][24] ) );
  DFFR_X1 \add_out_s2_reg[4][23]  ( .D(\add_out_s1[4][23] ), .CK(net18832), 
        .RN(RST), .Q(\add_out_s2[4][23] ) );
  DFFR_X1 \add_out_s2_reg[4][22]  ( .D(\add_out_s1[4][22] ), .CK(net18832), 
        .RN(RST), .Q(\add_out_s2[4][22] ) );
  DFFR_X1 \add_out_s2_reg[4][21]  ( .D(\add_out_s1[4][21] ), .CK(net18832), 
        .RN(RST), .Q(\add_out_s2[4][21] ) );
  DFFR_X1 \add_out_s2_reg[4][20]  ( .D(\add_out_s1[4][20] ), .CK(net18832), 
        .RN(RST), .Q(\add_out_s2[4][20] ) );
  DFFR_X1 \add_out_s2_reg[4][19]  ( .D(\add_out_s1[4][19] ), .CK(net18832), 
        .RN(RST), .Q(\add_out_s2[4][19] ) );
  DFFR_X1 \add_out_s2_reg[4][18]  ( .D(\add_out_s1[4][18] ), .CK(net18832), 
        .RN(RST), .Q(\add_out_s2[4][18] ) );
  DFFR_X1 \add_out_s2_reg[4][17]  ( .D(\add_out_s1[4][17] ), .CK(net18832), 
        .RN(RST), .Q(\add_out_s2[4][17] ) );
  DFFR_X1 \add_out_s2_reg[4][16]  ( .D(\add_out_s1[4][16] ), .CK(net18832), 
        .RN(RST), .Q(\add_out_s2[4][16] ) );
  DFFR_X1 \add_out_s2_reg[4][15]  ( .D(\add_out_s1[4][15] ), .CK(net18832), 
        .RN(RST), .Q(\add_out_s2[4][15] ) );
  DFFR_X1 \add_out_s2_reg[4][14]  ( .D(\add_out_s1[4][14] ), .CK(net18832), 
        .RN(RST), .Q(\add_out_s2[4][14] ) );
  DFFR_X1 \add_out_s2_reg[4][13]  ( .D(\add_out_s1[4][13] ), .CK(net18832), 
        .RN(RST), .Q(\add_out_s2[4][13] ) );
  DFFR_X1 \add_out_s2_reg[4][12]  ( .D(\add_out_s1[4][12] ), .CK(net18832), 
        .RN(RST), .Q(\add_out_s2[4][12] ) );
  DFFR_X1 \add_out_s2_reg[4][11]  ( .D(\add_out_s1[4][11] ), .CK(net18832), 
        .RN(RST), .Q(\add_out_s2[4][11] ) );
  DFFR_X1 \add_out_s2_reg[4][10]  ( .D(\add_out_s1[4][10] ), .CK(net18832), 
        .RN(RST), .Q(\add_out_s2[4][10] ) );
  DFFR_X1 \add_out_s2_reg[4][9]  ( .D(\add_out_s1[4][9] ), .CK(net18832), .RN(
        RST), .Q(\add_out_s2[4][9] ) );
  DFFR_X1 \add_out_s2_reg[4][8]  ( .D(\add_out_s1[4][8] ), .CK(net18832), .RN(
        RST), .Q(\add_out_s2[4][8] ) );
  DFFR_X1 \add_out_s2_reg[4][7]  ( .D(\add_out_s1[4][7] ), .CK(net18832), .RN(
        RST), .Q(\add_out_s2[4][7] ) );
  DFFR_X1 \add_out_s2_reg[4][6]  ( .D(\add_out_s1[4][6] ), .CK(net18832), .RN(
        RST), .Q(\add_out_s2[4][6] ) );
  DFFR_X1 \add_out_s2_reg[4][5]  ( .D(\add_out_s1[4][5] ), .CK(net18832), .RN(
        RST), .Q(\add_out_s2[4][5] ) );
  DFFR_X1 \add_out_s2_reg[4][4]  ( .D(\add_out_s1[4][4] ), .CK(net18832), .RN(
        RST), .Q(\add_out_s2[4][4] ) );
  DFFR_X1 \add_out_s2_reg[4][3]  ( .D(\add_out_s1[4][3] ), .CK(net18832), .RN(
        RST), .Q(\add_out_s2[4][3] ) );
  DFFR_X1 \add_out_s2_reg[4][2]  ( .D(\add_out_s1[4][2] ), .CK(net18832), .RN(
        RST), .Q(\add_out_s2[4][2] ) );
  DFFR_X1 \add_out_s2_reg[4][1]  ( .D(\add_out_s1[4][1] ), .CK(net18832), .RN(
        RST), .Q(\add_out_s2[4][1] ) );
  DFFR_X1 \add_out_s2_reg[4][0]  ( .D(\add_out_s1[4][0] ), .CK(net18832), .RN(
        RST), .Q(\add_out_s2[4][0] ) );
  DFFR_X1 \add_out_s3_reg[8][31]  ( .D(\add_out_s2[8][31] ), .CK(net18842), 
        .RN(RST), .Q(\add_out_s3[8][31] ) );
  DFFR_X1 \add_out_s3_reg[8][30]  ( .D(\add_out_s2[8][30] ), .CK(net18842), 
        .RN(RST), .Q(\add_out_s3[8][30] ) );
  DFFR_X1 \add_out_s3_reg[8][29]  ( .D(\add_out_s2[8][29] ), .CK(net18842), 
        .RN(RST), .Q(\add_out_s3[8][29] ) );
  DFFR_X1 \add_out_s3_reg[8][28]  ( .D(\add_out_s2[8][28] ), .CK(net18842), 
        .RN(RST), .Q(\add_out_s3[8][28] ) );
  DFFR_X1 \add_out_s3_reg[8][27]  ( .D(\add_out_s2[8][27] ), .CK(net18842), 
        .RN(RST), .Q(\add_out_s3[8][27] ) );
  DFFR_X1 \add_out_s3_reg[8][26]  ( .D(\add_out_s2[8][26] ), .CK(net18842), 
        .RN(RST), .Q(\add_out_s3[8][26] ) );
  DFFR_X1 \add_out_s3_reg[8][25]  ( .D(\add_out_s2[8][25] ), .CK(net18842), 
        .RN(RST), .Q(\add_out_s3[8][25] ) );
  DFFR_X1 \add_out_s3_reg[8][24]  ( .D(\add_out_s2[8][24] ), .CK(net18842), 
        .RN(RST), .Q(\add_out_s3[8][24] ) );
  DFFR_X1 \add_out_s3_reg[8][23]  ( .D(\add_out_s2[8][23] ), .CK(net18842), 
        .RN(RST), .Q(\add_out_s3[8][23] ) );
  DFFR_X1 \add_out_s3_reg[8][22]  ( .D(\add_out_s2[8][22] ), .CK(net18842), 
        .RN(RST), .Q(\add_out_s3[8][22] ) );
  DFFR_X1 \add_out_s3_reg[8][21]  ( .D(\add_out_s2[8][21] ), .CK(net18842), 
        .RN(RST), .Q(\add_out_s3[8][21] ) );
  DFFR_X1 \add_out_s3_reg[8][20]  ( .D(\add_out_s2[8][20] ), .CK(net18842), 
        .RN(RST), .Q(\add_out_s3[8][20] ) );
  DFFR_X1 \add_out_s3_reg[8][19]  ( .D(\add_out_s2[8][19] ), .CK(net18842), 
        .RN(RST), .Q(\add_out_s3[8][19] ) );
  DFFR_X1 \add_out_s3_reg[8][18]  ( .D(\add_out_s2[8][18] ), .CK(net18842), 
        .RN(RST), .Q(\add_out_s3[8][18] ) );
  DFFR_X1 \add_out_s3_reg[8][17]  ( .D(\add_out_s2[8][17] ), .CK(net18842), 
        .RN(RST), .Q(\add_out_s3[8][17] ) );
  DFFR_X1 \add_out_s3_reg[8][16]  ( .D(\add_out_s2[8][16] ), .CK(net18842), 
        .RN(RST), .Q(\add_out_s3[8][16] ) );
  DFFR_X1 \add_out_s3_reg[8][15]  ( .D(\add_out_s2[8][15] ), .CK(net18842), 
        .RN(RST), .Q(\add_out_s3[8][15] ) );
  DFFR_X1 \add_out_s3_reg[8][14]  ( .D(\add_out_s2[8][14] ), .CK(net18842), 
        .RN(RST), .Q(\add_out_s3[8][14] ) );
  DFFR_X1 \add_out_s3_reg[8][13]  ( .D(\add_out_s2[8][13] ), .CK(net18842), 
        .RN(RST), .Q(\add_out_s3[8][13] ) );
  DFFR_X1 \add_out_s3_reg[8][12]  ( .D(\add_out_s2[8][12] ), .CK(net18842), 
        .RN(RST), .Q(\add_out_s3[8][12] ) );
  DFFR_X1 \add_out_s3_reg[8][11]  ( .D(\add_out_s2[8][11] ), .CK(net18842), 
        .RN(RST), .Q(\add_out_s3[8][11] ) );
  DFFR_X1 \add_out_s3_reg[8][10]  ( .D(\add_out_s2[8][10] ), .CK(net18842), 
        .RN(RST), .Q(\add_out_s3[8][10] ) );
  DFFR_X1 \add_out_s3_reg[8][9]  ( .D(\add_out_s2[8][9] ), .CK(net18842), .RN(
        RST), .Q(\add_out_s3[8][9] ) );
  DFFR_X1 \add_out_s3_reg[8][8]  ( .D(\add_out_s2[8][8] ), .CK(net18842), .RN(
        RST), .Q(\add_out_s3[8][8] ) );
  DFFR_X1 \add_out_s3_reg[8][7]  ( .D(\add_out_s2[8][7] ), .CK(net18842), .RN(
        RST), .Q(\add_out_s3[8][7] ) );
  DFFR_X1 \add_out_s3_reg[8][6]  ( .D(\add_out_s2[8][6] ), .CK(net18842), .RN(
        RST), .Q(\add_out_s3[8][6] ) );
  DFFR_X1 \add_out_s3_reg[8][5]  ( .D(\add_out_s2[8][5] ), .CK(net18842), .RN(
        RST), .Q(\add_out_s3[8][5] ) );
  DFFR_X1 \add_out_s3_reg[8][4]  ( .D(\add_out_s2[8][4] ), .CK(net18842), .RN(
        RST), .Q(\add_out_s3[8][4] ) );
  DFFR_X1 \add_out_s3_reg[8][3]  ( .D(\add_out_s2[8][3] ), .CK(net18842), .RN(
        RST), .Q(\add_out_s3[8][3] ) );
  DFFR_X1 \add_out_s3_reg[8][2]  ( .D(\add_out_s2[8][2] ), .CK(net18842), .RN(
        RST), .Q(\add_out_s3[8][2] ) );
  DFFR_X1 \add_out_s3_reg[8][1]  ( .D(\add_out_s2[8][1] ), .CK(net18842), .RN(
        RST), .Q(\add_out_s3[8][1] ) );
  DFFR_X1 \add_out_s3_reg[8][0]  ( .D(\add_out_s2[8][0] ), .CK(net18842), .RN(
        RST), .Q(\add_out_s3[8][0] ) );
  DFFR_X1 \add_out_s4_reg[12][0]  ( .D(\add_out_s3[12][0] ), .CK(net18822), 
        .RN(RST), .Q(\add_out_s4[12][0] ) );
  DFFR_X1 \add_out_s4_reg[12][1]  ( .D(\add_out_s3[12][1] ), .CK(net18822), 
        .RN(RST), .Q(\add_out_s4[12][1] ) );
  DFFR_X1 \add_out_s4_reg[12][2]  ( .D(\add_out_s3[12][2] ), .CK(net18822), 
        .RN(RST), .Q(\add_out_s4[12][2] ) );
  DFFR_X1 \add_out_s4_reg[12][3]  ( .D(\add_out_s3[12][3] ), .CK(net18822), 
        .RN(RST), .Q(\add_out_s4[12][3] ) );
  DFFR_X1 \add_out_s4_reg[12][4]  ( .D(\add_out_s3[12][4] ), .CK(net18822), 
        .RN(RST), .Q(\add_out_s4[12][4] ) );
  DFFR_X1 \add_out_s4_reg[12][5]  ( .D(\add_out_s3[12][5] ), .CK(net18822), 
        .RN(RST), .Q(\add_out_s4[12][5] ) );
  DFFR_X1 \add_out_s4_reg[12][6]  ( .D(\add_out_s3[12][6] ), .CK(net18822), 
        .RN(RST), .Q(\add_out_s4[12][6] ) );
  DFFR_X1 \add_out_s4_reg[12][7]  ( .D(\add_out_s3[12][7] ), .CK(net18822), 
        .RN(RST), .Q(\add_out_s4[12][7] ) );
  DFFR_X1 \add_out_s4_reg[12][8]  ( .D(\add_out_s3[12][8] ), .CK(net18822), 
        .RN(RST), .Q(\add_out_s4[12][8] ) );
  DFFR_X1 \add_out_s4_reg[12][9]  ( .D(\add_out_s3[12][9] ), .CK(net18822), 
        .RN(RST), .Q(\add_out_s4[12][9] ) );
  DFFR_X1 \add_out_s4_reg[12][10]  ( .D(\add_out_s3[12][10] ), .CK(net18822), 
        .RN(RST), .Q(\add_out_s4[12][10] ) );
  DFFR_X1 \add_out_s4_reg[12][11]  ( .D(\add_out_s3[12][11] ), .CK(net18822), 
        .RN(RST), .Q(\add_out_s4[12][11] ) );
  DFFR_X1 \add_out_s4_reg[12][12]  ( .D(\add_out_s3[12][12] ), .CK(net18822), 
        .RN(RST), .Q(\add_out_s4[12][12] ) );
  DFFR_X1 \add_out_s4_reg[12][13]  ( .D(\add_out_s3[12][13] ), .CK(net18822), 
        .RN(RST), .Q(\add_out_s4[12][13] ) );
  DFFR_X1 \add_out_s4_reg[12][14]  ( .D(\add_out_s3[12][14] ), .CK(net18822), 
        .RN(RST), .Q(\add_out_s4[12][14] ) );
  DFFR_X1 \add_out_s4_reg[12][15]  ( .D(\add_out_s3[12][15] ), .CK(net18822), 
        .RN(RST), .Q(\add_out_s4[12][15] ) );
  DFFR_X1 \add_out_s4_reg[12][16]  ( .D(\add_out_s3[12][16] ), .CK(net18822), 
        .RN(RST), .Q(\add_out_s4[12][16] ) );
  DFFR_X1 \add_out_s4_reg[12][17]  ( .D(\add_out_s3[12][17] ), .CK(net18822), 
        .RN(RST), .Q(\add_out_s4[12][17] ) );
  DFFR_X1 \add_out_s4_reg[12][18]  ( .D(\add_out_s3[12][18] ), .CK(net18822), 
        .RN(RST), .Q(\add_out_s4[12][18] ) );
  DFFR_X1 \add_out_s4_reg[12][19]  ( .D(\add_out_s3[12][19] ), .CK(net18822), 
        .RN(RST), .Q(\add_out_s4[12][19] ) );
  DFFR_X1 \add_out_s4_reg[12][20]  ( .D(\add_out_s3[12][20] ), .CK(net18822), 
        .RN(RST), .Q(\add_out_s4[12][20] ) );
  DFFR_X1 \add_out_s4_reg[12][21]  ( .D(\add_out_s3[12][21] ), .CK(net18822), 
        .RN(RST), .Q(\add_out_s4[12][21] ) );
  DFFR_X1 \add_out_s4_reg[12][22]  ( .D(\add_out_s3[12][22] ), .CK(net18822), 
        .RN(RST), .Q(\add_out_s4[12][22] ) );
  DFFR_X1 \add_out_s4_reg[12][23]  ( .D(\add_out_s3[12][23] ), .CK(net18822), 
        .RN(RST), .Q(\add_out_s4[12][23] ) );
  DFFR_X1 \add_out_s4_reg[12][24]  ( .D(\add_out_s3[12][24] ), .CK(net18822), 
        .RN(RST), .Q(\add_out_s4[12][24] ) );
  DFFR_X1 \add_out_s4_reg[12][25]  ( .D(\add_out_s3[12][25] ), .CK(net18822), 
        .RN(RST), .Q(\add_out_s4[12][25] ) );
  DFFR_X1 \add_out_s4_reg[12][26]  ( .D(\add_out_s3[12][26] ), .CK(net18822), 
        .RN(RST), .Q(\add_out_s4[12][26] ) );
  DFFR_X1 \add_out_s4_reg[12][27]  ( .D(\add_out_s3[12][27] ), .CK(net18822), 
        .RN(RST), .Q(\add_out_s4[12][27] ) );
  DFFR_X1 \add_out_s4_reg[12][28]  ( .D(\add_out_s3[12][28] ), .CK(net18822), 
        .RN(RST), .Q(\add_out_s4[12][28] ) );
  DFFR_X1 \add_out_s4_reg[12][29]  ( .D(\add_out_s3[12][29] ), .CK(net18822), 
        .RN(RST), .Q(\add_out_s4[12][29] ) );
  DFFR_X1 \add_out_s4_reg[12][30]  ( .D(\add_out_s3[12][30] ), .CK(net18822), 
        .RN(RST), .Q(\add_out_s4[12][30] ) );
  DFFR_X1 \add_out_s4_reg[12][31]  ( .D(\add_out_s3[12][31] ), .CK(net18822), 
        .RN(RST), .Q(\add_out_s4[12][31] ) );
  HA_X1 \sub_x_1/U31  ( .A(n43), .B(n74), .CO(\sub_x_1/n29 ), .S(
        \A_shifted[-32][34] ) );
  HA_X1 \sub_x_1/U18  ( .A(\sub_x_1/n17 ), .B(n66), .CO(\sub_x_1/n16 ), .S(
        \A_shifted[-32][47] ) );
  HA_X1 \sub_x_1/U12  ( .A(\sub_x_1/n11 ), .B(n62), .CO(\sub_x_1/n10 ), .S(
        \A_shifted[-32][53] ) );
  HA_X1 \sub_x_1/U10  ( .A(\sub_x_1/n9 ), .B(n79), .CO(\sub_x_1/n8 ), .S(
        \A_shifted[-32][55] ) );
  HA_X1 \sub_x_1/U9  ( .A(\sub_x_1/n8 ), .B(n78), .CO(\sub_x_1/n7 ), .S(
        \A_shifted[-32][56] ) );
  HA_X1 \sub_x_1/U8  ( .A(\sub_x_1/n7 ), .B(n60), .CO(\sub_x_1/n6 ), .S(
        \A_shifted[-32][57] ) );
  HA_X1 \sub_x_1/U7  ( .A(\sub_x_1/n6 ), .B(n59), .CO(\sub_x_1/n5 ), .S(
        \A_shifted[-32][58] ) );
  HA_X1 \sub_x_1/U6  ( .A(\sub_x_1/n5 ), .B(n58), .CO(\sub_x_1/n4 ), .S(
        \A_shifted[-32][59] ) );
  DFFR_X1 \add_out_s2_reg[4][28]  ( .D(\add_out_s1[4][28] ), .CK(net18832), 
        .RN(RST), .Q(\add_out_s2[4][28] ) );
  DFFR_X1 \add_out_s2_reg[4][29]  ( .D(\add_out_s1[4][29] ), .CK(net18832), 
        .RN(RST), .Q(\add_out_s2[4][29] ) );
  DFFR_X1 \add_out_s2_reg[4][30]  ( .D(\add_out_s1[4][30] ), .CK(net18832), 
        .RN(RST), .Q(\add_out_s2[4][30] ) );
  DFFR_X1 \add_out_s2_reg[4][31]  ( .D(\add_out_s1[4][31] ), .CK(net18832), 
        .RN(RST), .Q(\add_out_s2[4][31] ) );
  DFFRS_X1 \add_out_s2_reg[4][27]  ( .D(\add_out_s1[4][27] ), .CK(net18832), 
        .RN(RST), .SN(1'b1), .Q(\add_out_s2[4][27] ) );
  NAND3_X1 U5 ( .A1(n65), .A2(n80), .A3(\sub_x_1/n16 ), .ZN(n2) );
  NOR2_X1 U6 ( .A1(\sub_x_1/B[21] ), .A2(n2), .ZN(\sub_x_1/n11 ) );
  XOR2_X1 U7 ( .A(\sub_x_1/B[21] ), .B(n2), .Z(\A_shifted[-32][52] ) );
  NAND3_X1 U8 ( .A1(\sub_x_1/n26 ), .A2(n87), .A3(n37), .ZN(n3) );
  XNOR2_X1 U9 ( .A(n3), .B(n68), .ZN(\A_shifted[-32][42] ) );
  XNOR2_X1 U10 ( .A(\sub_x_1/n4 ), .B(A[29]), .ZN(\A_shifted[-32][60] ) );
  INV_X1 U11 ( .A(\sub_x_1/n4 ), .ZN(n4) );
  NOR2_X1 U12 ( .A1(A[29]), .A2(n4), .ZN(\sub_x_1/n3 ) );
  NAND2_X1 U13 ( .A1(n64), .A2(\sub_x_1/n15 ), .ZN(n5) );
  XOR2_X1 U14 ( .A(A[19]), .B(n5), .Z(\A_shifted[-32][50] ) );
  NOR3_X1 U15 ( .A1(n89), .A2(n85), .A3(A[14]), .ZN(n6) );
  XNOR2_X1 U16 ( .A(\sub_x_1/B[15] ), .B(n6), .ZN(\A_shifted[-32][46] ) );
  XNOR2_X1 U17 ( .A(\sub_x_1/n3 ), .B(A[30]), .ZN(\A_shifted[-32][61] ) );
  INV_X1 U18 ( .A(\sub_x_1/n3 ), .ZN(n7) );
  NOR2_X1 U19 ( .A1(A[30]), .A2(n7), .ZN(\sub_x_1/n2 ) );
  NAND3_X1 U20 ( .A1(\sub_x_1/n15 ), .A2(n63), .A3(n64), .ZN(n8) );
  XOR2_X1 U21 ( .A(A[20]), .B(n8), .Z(\A_shifted[-32][51] ) );
  XOR2_X1 U22 ( .A(A[10]), .B(n89), .Z(\A_shifted[-32][41] ) );
  INV_X1 U23 ( .A(A[20]), .ZN(n9) );
  AND3_X1 U24 ( .A1(n64), .A2(n63), .A3(n9), .ZN(n80) );
  NAND2_X1 U25 ( .A1(n69), .A2(\sub_x_1/n25 ), .ZN(n10) );
  XOR2_X1 U26 ( .A(A[9]), .B(n10), .Z(\A_shifted[-32][40] ) );
  BUF_X4 U27 ( .A(A[2]), .Z(n625) );
  AND2_X1 U29 ( .A1(\sub_x_1/n17 ), .A2(n66), .ZN(n12) );
  BUF_X1 U30 ( .A(\A_shifted[-32][45] ), .Z(n52) );
  BUF_X1 U31 ( .A(\A_shifted[-32][36] ), .Z(n629) );
  BUF_X2 U32 ( .A(A[1]), .Z(n636) );
  BUF_X2 U33 ( .A(A[0]), .Z(n635) );
  BUF_X1 U34 ( .A(A[3]), .Z(n626) );
  BUF_X2 U35 ( .A(A[4]), .Z(n637) );
  BUF_X1 U36 ( .A(A[6]), .Z(n639) );
  BUF_X1 U37 ( .A(\A_shifted[-32][51] ), .Z(n33) );
  BUF_X1 U38 ( .A(\A_shifted[-32][46] ), .Z(n50) );
  BUF_X1 U39 ( .A(\A_shifted[-32][40] ), .Z(n54) );
  BUF_X1 U40 ( .A(\A_shifted[-32][47] ), .Z(n90) );
  BUF_X1 U41 ( .A(\A_shifted[-32][43] ), .Z(n55) );
  BUF_X1 U42 ( .A(\A_shifted[-32][38] ), .Z(n632) );
  BUF_X1 U43 ( .A(\A_shifted[-32][42] ), .Z(n96) );
  BUF_X1 U44 ( .A(\A_shifted[-32][36] ), .Z(n630) );
  AND2_X1 U45 ( .A1(n49), .A2(n70), .ZN(\sub_x_1/n25 ) );
  XNOR2_X1 U46 ( .A(n47), .B(A[5]), .ZN(\A_shifted[-32][36] ) );
  AND2_X1 U47 ( .A1(n48), .A2(n71), .ZN(\sub_x_1/n26 ) );
  BUF_X2 U48 ( .A(\A_shifted[-32][37] ), .Z(n17) );
  BUF_X2 U49 ( .A(\A_shifted[-32][34] ), .Z(n23) );
  NOR2_X1 U50 ( .A1(A[9]), .A2(A[8]), .ZN(n36) );
  BUF_X2 U51 ( .A(\A_shifted[-32][33] ), .Z(n18) );
  BUF_X2 U52 ( .A(\A_shifted[-32][35] ), .Z(n19) );
  AND3_X1 U53 ( .A1(n45), .A2(n73), .A3(n72), .ZN(n48) );
  AND2_X1 U54 ( .A1(n71), .A2(n72), .ZN(n34) );
  CLKBUF_X1 U55 ( .A(A[5]), .Z(n638) );
  CLKBUF_X1 U56 ( .A(A[7]), .Z(n640) );
  INV_X1 U57 ( .A(A[2]), .ZN(n75) );
  BUF_X1 U58 ( .A(\A_shifted[-32][54] ), .Z(n57) );
  BUF_X1 U59 ( .A(\A_shifted[-32][53] ), .Z(n32) );
  BUF_X1 U60 ( .A(\A_shifted[-32][50] ), .Z(n95) );
  BUF_X1 U61 ( .A(\A_shifted[-32][49] ), .Z(n41) );
  BUF_X1 U62 ( .A(\A_shifted[-32][52] ), .Z(n53) );
  BUF_X1 U63 ( .A(\A_shifted[-32][41] ), .Z(n94) );
  BUF_X1 U64 ( .A(\A_shifted[-32][48] ), .Z(n93) );
  BUF_X1 U65 ( .A(\A_shifted[-32][44] ), .Z(n92) );
  BUF_X1 U66 ( .A(\A_shifted[-32][44] ), .Z(n91) );
  BUF_X1 U67 ( .A(\A_shifted[-32][39] ), .Z(n634) );
  XNOR2_X1 U68 ( .A(\sub_x_1/n21 ), .B(A[12]), .ZN(\A_shifted[-32][43] ) );
  XNOR2_X1 U69 ( .A(n49), .B(A[7]), .ZN(\A_shifted[-32][38] ) );
  AND2_X1 U70 ( .A1(\sub_x_1/n26 ), .A2(n70), .ZN(n51) );
  XNOR2_X1 U71 ( .A(n48), .B(A[6]), .ZN(\A_shifted[-32][37] ) );
  AND2_X1 U72 ( .A1(n37), .A2(n88), .ZN(n35) );
  BUF_X1 U73 ( .A(B[25]), .Z(n44) );
  OR2_X1 U74 ( .A1(n39), .A2(A[12]), .ZN(n38) );
  BUF_X1 U75 ( .A(B[9]), .Z(n46) );
  XNOR2_X1 U76 ( .A(A[4]), .B(n45), .ZN(\A_shifted[-32][35] ) );
  XNOR2_X1 U77 ( .A(n625), .B(n42), .ZN(\A_shifted[-32][33] ) );
  XNOR2_X1 U78 ( .A(n635), .B(n76), .ZN(\A_shifted[-32][32] ) );
  NAND2_X1 U79 ( .A1(n68), .A2(n82), .ZN(n39) );
  AND2_X1 U80 ( .A1(n69), .A2(n70), .ZN(n37) );
  AND3_X1 U81 ( .A1(n42), .A2(n75), .A3(n74), .ZN(n45) );
  BUF_X1 U82 ( .A(A[22]), .Z(\sub_x_1/B[22] ) );
  BUF_X1 U83 ( .A(A[21]), .Z(\sub_x_1/B[21] ) );
  NOR2_X1 U84 ( .A1(A[1]), .A2(A[0]), .ZN(n42) );
  BUF_X1 U85 ( .A(A[10]), .Z(n642) );
  BUF_X1 U86 ( .A(A[17]), .Z(\sub_x_1/B[17] ) );
  INV_X1 U87 ( .A(A[1]), .ZN(n76) );
  BUF_X1 U88 ( .A(A[3]), .Z(n627) );
  BUF_X1 U89 ( .A(A[8]), .Z(n641) );
  BUF_X1 U90 ( .A(A[11]), .Z(n643) );
  AND2_X1 U91 ( .A1(n29), .A2(n77), .ZN(n43) );
  NOR2_X1 U92 ( .A1(A[2]), .A2(A[1]), .ZN(n29) );
  AND2_X1 U93 ( .A1(n47), .A2(n34), .ZN(n49) );
  NOR2_X1 U94 ( .A1(n38), .A2(n30), .ZN(n40) );
  NAND2_X1 U95 ( .A1(n31), .A2(n87), .ZN(n30) );
  NOR2_X1 U96 ( .A1(A[14]), .A2(\sub_x_1/B[15] ), .ZN(n31) );
  AND2_X1 U97 ( .A1(\sub_x_1/n26 ), .A2(n35), .ZN(\sub_x_1/n21 ) );
  AND2_X1 U98 ( .A1(\sub_x_1/n26 ), .A2(n37), .ZN(\sub_x_1/n24 ) );
  NAND2_X1 U99 ( .A1(\sub_x_1/n25 ), .A2(n36), .ZN(n89) );
  XNOR2_X1 U100 ( .A(n51), .B(A[8]), .ZN(\A_shifted[-32][39] ) );
  AND2_X1 U101 ( .A1(\sub_x_1/n24 ), .A2(n40), .ZN(\sub_x_1/n17 ) );
  AND2_X1 U102 ( .A1(n12), .A2(n65), .ZN(\sub_x_1/n15 ) );
  XNOR2_X1 U103 ( .A(\sub_x_1/n15 ), .B(A[18]), .ZN(\A_shifted[-32][49] ) );
  AND2_X1 U104 ( .A1(\sub_x_1/n29 ), .A2(n73), .ZN(n47) );
  XNOR2_X1 U105 ( .A(\sub_x_1/n19 ), .B(A[14]), .ZN(\A_shifted[-32][45] ) );
  XOR2_X1 U106 ( .A(\sub_x_1/n6 ), .B(n59), .Z(n56) );
  XNOR2_X1 U107 ( .A(\sub_x_1/n10 ), .B(\sub_x_1/B[23] ), .ZN(
        \A_shifted[-32][54] ) );
  XNOR2_X1 U108 ( .A(A[31]), .B(\sub_x_1/n2 ), .ZN(\A_shifted[-32][62] ) );
  INV_X1 U109 ( .A(A[28]), .ZN(n58) );
  INV_X1 U110 ( .A(A[27]), .ZN(n59) );
  INV_X1 U111 ( .A(A[26]), .ZN(n60) );
  INV_X1 U112 ( .A(\sub_x_1/B[23] ), .ZN(n61) );
  INV_X1 U113 ( .A(\sub_x_1/B[22] ), .ZN(n62) );
  INV_X1 U114 ( .A(A[19]), .ZN(n63) );
  INV_X1 U115 ( .A(A[18]), .ZN(n64) );
  INV_X1 U116 ( .A(\sub_x_1/B[17] ), .ZN(n65) );
  INV_X1 U117 ( .A(A[16]), .ZN(n66) );
  INV_X1 U118 ( .A(A[12]), .ZN(n67) );
  INV_X1 U119 ( .A(A[11]), .ZN(n68) );
  INV_X1 U120 ( .A(A[8]), .ZN(n69) );
  INV_X1 U121 ( .A(A[0]), .ZN(n77) );
  INV_X1 U122 ( .A(A[25]), .ZN(n78) );
  INV_X1 U123 ( .A(A[24]), .ZN(n79) );
  NOR2_X1 U124 ( .A1(n89), .A2(n85), .ZN(\sub_x_1/n19 ) );
  NAND2_X1 U125 ( .A1(\sub_x_1/n21 ), .A2(n67), .ZN(n81) );
  INV_X1 U126 ( .A(A[13]), .ZN(n82) );
  NOR2_X1 U127 ( .A1(A[10]), .A2(A[9]), .ZN(n87) );
  NOR2_X1 U128 ( .A1(A[10]), .A2(A[11]), .ZN(n84) );
  NOR2_X1 U129 ( .A1(A[13]), .A2(A[12]), .ZN(n83) );
  NAND2_X1 U130 ( .A1(n84), .A2(n83), .ZN(n85) );
  INV_X1 U131 ( .A(n84), .ZN(n86) );
  NOR2_X1 U132 ( .A1(n86), .A2(A[9]), .ZN(n88) );
  INV_X1 U133 ( .A(A[7]), .ZN(n70) );
  INV_X1 U134 ( .A(A[5]), .ZN(n72) );
  INV_X1 U135 ( .A(A[6]), .ZN(n71) );
  AND2_X1 U136 ( .A1(\sub_x_1/n10 ), .A2(n61), .ZN(\sub_x_1/n9 ) );
  INV_X1 U137 ( .A(A[3]), .ZN(n74) );
  XNOR2_X1 U138 ( .A(n12), .B(\sub_x_1/B[17] ), .ZN(\A_shifted[-32][48] ) );
  INV_X1 U139 ( .A(A[4]), .ZN(n73) );
  XNOR2_X1 U140 ( .A(n81), .B(n82), .ZN(\A_shifted[-32][44] ) );
  BUF_X2 U141 ( .A(\A_shifted[-32][32] ), .Z(n628) );
  BUF_X2 U142 ( .A(\A_shifted[-32][38] ), .Z(n631) );
  BUF_X2 U143 ( .A(\A_shifted[-32][39] ), .Z(n633) );
  BUF_X2 U144 ( .A(A[15]), .Z(\sub_x_1/B[15] ) );
  BUF_X1 U145 ( .A(A[23]), .Z(\sub_x_1/B[23] ) );
endmodule


module MUX_2to1_N32_5 ( IN0, IN1, SEL, Y );
  input [31:0] IN0;
  input [31:0] IN1;
  output [31:0] Y;
  input SEL;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12;

  MUX2_X1 U1 ( .A(IN0[10]), .B(IN1[10]), .S(n9), .Z(Y[10]) );
  MUX2_X1 U2 ( .A(IN0[9]), .B(IN1[9]), .S(n9), .Z(Y[9]) );
  MUX2_X1 U3 ( .A(IN0[13]), .B(IN1[13]), .S(SEL), .Z(Y[13]) );
  MUX2_X1 U4 ( .A(IN0[30]), .B(IN1[30]), .S(n9), .Z(Y[30]) );
  MUX2_X1 U5 ( .A(IN0[18]), .B(IN1[18]), .S(SEL), .Z(Y[18]) );
  MUX2_X1 U6 ( .A(IN0[7]), .B(IN1[7]), .S(n9), .Z(Y[7]) );
  MUX2_X2 U7 ( .A(IN0[11]), .B(IN1[11]), .S(SEL), .Z(Y[11]) );
  INV_X1 U8 ( .A(n10), .ZN(n9) );
  INV_X1 U9 ( .A(SEL), .ZN(n10) );
  NAND2_X1 U10 ( .A1(n2), .A2(n1), .ZN(Y[28]) );
  NAND2_X1 U11 ( .A1(IN1[28]), .A2(n9), .ZN(n1) );
  NAND2_X1 U12 ( .A1(IN0[28]), .A2(n10), .ZN(n2) );
  NAND2_X1 U13 ( .A1(n4), .A2(n3), .ZN(Y[24]) );
  NAND2_X1 U14 ( .A1(IN1[24]), .A2(SEL), .ZN(n3) );
  NAND2_X1 U15 ( .A1(IN0[24]), .A2(n10), .ZN(n4) );
  NAND2_X1 U16 ( .A1(n6), .A2(n5), .ZN(Y[25]) );
  NAND2_X1 U17 ( .A1(n9), .A2(IN1[25]), .ZN(n5) );
  NAND2_X1 U18 ( .A1(IN0[25]), .A2(n10), .ZN(n6) );
  NAND2_X1 U19 ( .A1(n8), .A2(n7), .ZN(Y[31]) );
  NAND2_X1 U20 ( .A1(IN0[31]), .A2(n10), .ZN(n7) );
  NAND2_X1 U21 ( .A1(IN1[31]), .A2(n9), .ZN(n8) );
  NAND2_X1 U22 ( .A1(n12), .A2(n11), .ZN(Y[0]) );
  NAND2_X1 U23 ( .A1(IN1[0]), .A2(SEL), .ZN(n11) );
  NAND2_X1 U24 ( .A1(IN0[0]), .A2(n10), .ZN(n12) );
  MUX2_X1 U25 ( .A(IN0[12]), .B(IN1[12]), .S(SEL), .Z(Y[12]) );
  MUX2_X1 U26 ( .A(IN0[14]), .B(IN1[14]), .S(SEL), .Z(Y[14]) );
  MUX2_X1 U27 ( .A(IN0[15]), .B(IN1[15]), .S(SEL), .Z(Y[15]) );
  MUX2_X1 U28 ( .A(IN0[16]), .B(IN1[16]), .S(SEL), .Z(Y[16]) );
  MUX2_X1 U29 ( .A(IN0[17]), .B(IN1[17]), .S(SEL), .Z(Y[17]) );
  MUX2_X1 U30 ( .A(IN0[19]), .B(IN1[19]), .S(SEL), .Z(Y[19]) );
  MUX2_X1 U31 ( .A(IN0[1]), .B(IN1[1]), .S(SEL), .Z(Y[1]) );
  MUX2_X1 U32 ( .A(IN0[20]), .B(IN1[20]), .S(SEL), .Z(Y[20]) );
  MUX2_X1 U33 ( .A(IN0[21]), .B(IN1[21]), .S(SEL), .Z(Y[21]) );
  MUX2_X1 U34 ( .A(IN0[22]), .B(IN1[22]), .S(SEL), .Z(Y[22]) );
  MUX2_X1 U35 ( .A(IN0[23]), .B(IN1[23]), .S(SEL), .Z(Y[23]) );
  MUX2_X1 U36 ( .A(IN0[26]), .B(IN1[26]), .S(n9), .Z(Y[26]) );
  MUX2_X1 U37 ( .A(IN0[27]), .B(IN1[27]), .S(n9), .Z(Y[27]) );
  MUX2_X1 U38 ( .A(IN0[29]), .B(IN1[29]), .S(n9), .Z(Y[29]) );
  MUX2_X1 U39 ( .A(IN0[2]), .B(IN1[2]), .S(n9), .Z(Y[2]) );
  MUX2_X1 U40 ( .A(IN0[3]), .B(IN1[3]), .S(n9), .Z(Y[3]) );
  MUX2_X1 U41 ( .A(IN0[4]), .B(IN1[4]), .S(n9), .Z(Y[4]) );
  MUX2_X1 U42 ( .A(IN0[5]), .B(IN1[5]), .S(n9), .Z(Y[5]) );
  MUX2_X1 U43 ( .A(IN0[6]), .B(IN1[6]), .S(n9), .Z(Y[6]) );
  MUX2_X1 U44 ( .A(IN0[8]), .B(IN1[8]), .S(n9), .Z(Y[8]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_reg_N32_6 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18782, net18784, net18786, net18787, net18790, net18793;
  assign net18782 = EN;
  assign net18784 = CLK;
  assign ENCLK = net18786;
  assign net18793 = TE;

  DLL_X1 latch ( .D(net18787), .GN(net18784), .Q(net18790) );
  AND2_X1 main_gate ( .A1(net18790), .A2(net18784), .ZN(net18786) );
  OR2_X1 test_or ( .A1(net18782), .A2(net18793), .ZN(net18787) );
endmodule


module reg_N32_6 ( D, Q, EN, CLK, RST );
  input [31:0] D;
  output [31:0] Q;
  input EN, CLK, RST;
  wire   net18798;

  SNPS_CLOCK_GATE_HIGH_reg_N32_6 clk_gate_Q_reg ( .CLK(CLK), .EN(EN), .ENCLK(
        net18798), .TE(1'b0) );
  DFFR_X1 \Q_reg[31]  ( .D(D[31]), .CK(net18798), .RN(RST), .Q(Q[31]) );
  DFFR_X1 \Q_reg[30]  ( .D(D[30]), .CK(net18798), .RN(RST), .Q(Q[30]) );
  DFFR_X1 \Q_reg[29]  ( .D(D[29]), .CK(net18798), .RN(RST), .Q(Q[29]) );
  DFFR_X1 \Q_reg[28]  ( .D(D[28]), .CK(net18798), .RN(RST), .Q(Q[28]) );
  DFFR_X1 \Q_reg[27]  ( .D(D[27]), .CK(net18798), .RN(RST), .Q(Q[27]) );
  DFFR_X1 \Q_reg[26]  ( .D(D[26]), .CK(net18798), .RN(RST), .Q(Q[26]) );
  DFFR_X1 \Q_reg[25]  ( .D(D[25]), .CK(net18798), .RN(RST), .Q(Q[25]) );
  DFFR_X1 \Q_reg[24]  ( .D(D[24]), .CK(net18798), .RN(RST), .Q(Q[24]) );
  DFFR_X1 \Q_reg[23]  ( .D(D[23]), .CK(net18798), .RN(RST), .Q(Q[23]) );
  DFFR_X1 \Q_reg[22]  ( .D(D[22]), .CK(net18798), .RN(RST), .Q(Q[22]) );
  DFFR_X1 \Q_reg[21]  ( .D(D[21]), .CK(net18798), .RN(RST), .Q(Q[21]) );
  DFFR_X1 \Q_reg[20]  ( .D(D[20]), .CK(net18798), .RN(RST), .Q(Q[20]) );
  DFFR_X1 \Q_reg[19]  ( .D(D[19]), .CK(net18798), .RN(RST), .Q(Q[19]) );
  DFFR_X1 \Q_reg[18]  ( .D(D[18]), .CK(net18798), .RN(RST), .Q(Q[18]) );
  DFFR_X1 \Q_reg[17]  ( .D(D[17]), .CK(net18798), .RN(RST), .Q(Q[17]) );
  DFFR_X1 \Q_reg[16]  ( .D(D[16]), .CK(net18798), .RN(RST), .Q(Q[16]) );
  DFFR_X1 \Q_reg[15]  ( .D(D[15]), .CK(net18798), .RN(RST), .Q(Q[15]) );
  DFFR_X1 \Q_reg[14]  ( .D(D[14]), .CK(net18798), .RN(RST), .Q(Q[14]) );
  DFFR_X1 \Q_reg[13]  ( .D(D[13]), .CK(net18798), .RN(RST), .Q(Q[13]) );
  DFFR_X1 \Q_reg[12]  ( .D(D[12]), .CK(net18798), .RN(RST), .Q(Q[12]) );
  DFFR_X1 \Q_reg[11]  ( .D(D[11]), .CK(net18798), .RN(RST), .Q(Q[11]) );
  DFFR_X1 \Q_reg[10]  ( .D(D[10]), .CK(net18798), .RN(RST), .Q(Q[10]) );
  DFFR_X1 \Q_reg[9]  ( .D(D[9]), .CK(net18798), .RN(RST), .Q(Q[9]) );
  DFFR_X1 \Q_reg[8]  ( .D(D[8]), .CK(net18798), .RN(RST), .Q(Q[8]) );
  DFFR_X1 \Q_reg[7]  ( .D(D[7]), .CK(net18798), .RN(RST), .Q(Q[7]) );
  DFFR_X1 \Q_reg[6]  ( .D(D[6]), .CK(net18798), .RN(RST), .Q(Q[6]) );
  DFFR_X1 \Q_reg[5]  ( .D(D[5]), .CK(net18798), .RN(RST), .Q(Q[5]) );
  DFFR_X1 \Q_reg[4]  ( .D(D[4]), .CK(net18798), .RN(RST), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(D[3]), .CK(net18798), .RN(RST), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(D[2]), .CK(net18798), .RN(RST), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(D[1]), .CK(net18798), .RN(RST), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(D[0]), .CK(net18798), .RN(RST), .Q(Q[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_reg_N32_5 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18782, net18784, net18786, net18787, net18790, net18793;
  assign net18782 = EN;
  assign net18784 = CLK;
  assign ENCLK = net18786;
  assign net18793 = TE;

  DLL_X1 latch ( .D(net18787), .GN(net18784), .Q(net18790) );
  AND2_X1 main_gate ( .A1(net18790), .A2(net18784), .ZN(net18786) );
  OR2_X1 test_or ( .A1(net18782), .A2(net18793), .ZN(net18787) );
endmodule


module reg_N32_5 ( D, Q, EN, CLK, RST );
  input [31:0] D;
  output [31:0] Q;
  input EN, CLK, RST;
  wire   net18798;

  SNPS_CLOCK_GATE_HIGH_reg_N32_5 clk_gate_Q_reg ( .CLK(CLK), .EN(EN), .ENCLK(
        net18798), .TE(1'b0) );
  DFFR_X1 \Q_reg[31]  ( .D(D[31]), .CK(net18798), .RN(RST), .Q(Q[31]) );
  DFFR_X1 \Q_reg[30]  ( .D(D[30]), .CK(net18798), .RN(RST), .Q(Q[30]) );
  DFFR_X1 \Q_reg[29]  ( .D(D[29]), .CK(net18798), .RN(RST), .Q(Q[29]) );
  DFFR_X1 \Q_reg[28]  ( .D(D[28]), .CK(net18798), .RN(RST), .Q(Q[28]) );
  DFFR_X1 \Q_reg[27]  ( .D(D[27]), .CK(net18798), .RN(RST), .Q(Q[27]) );
  DFFR_X1 \Q_reg[26]  ( .D(D[26]), .CK(net18798), .RN(RST), .Q(Q[26]) );
  DFFR_X1 \Q_reg[25]  ( .D(D[25]), .CK(net18798), .RN(RST), .Q(Q[25]) );
  DFFR_X1 \Q_reg[24]  ( .D(D[24]), .CK(net18798), .RN(RST), .Q(Q[24]) );
  DFFR_X1 \Q_reg[23]  ( .D(D[23]), .CK(net18798), .RN(RST), .Q(Q[23]) );
  DFFR_X1 \Q_reg[22]  ( .D(D[22]), .CK(net18798), .RN(RST), .Q(Q[22]) );
  DFFR_X1 \Q_reg[21]  ( .D(D[21]), .CK(net18798), .RN(RST), .Q(Q[21]) );
  DFFR_X1 \Q_reg[20]  ( .D(D[20]), .CK(net18798), .RN(RST), .Q(Q[20]) );
  DFFR_X1 \Q_reg[19]  ( .D(D[19]), .CK(net18798), .RN(RST), .Q(Q[19]) );
  DFFR_X1 \Q_reg[18]  ( .D(D[18]), .CK(net18798), .RN(RST), .Q(Q[18]) );
  DFFR_X1 \Q_reg[17]  ( .D(D[17]), .CK(net18798), .RN(RST), .Q(Q[17]) );
  DFFR_X1 \Q_reg[16]  ( .D(D[16]), .CK(net18798), .RN(RST), .Q(Q[16]) );
  DFFR_X1 \Q_reg[15]  ( .D(D[15]), .CK(net18798), .RN(RST), .Q(Q[15]) );
  DFFR_X1 \Q_reg[14]  ( .D(D[14]), .CK(net18798), .RN(RST), .Q(Q[14]) );
  DFFR_X1 \Q_reg[13]  ( .D(D[13]), .CK(net18798), .RN(RST), .Q(Q[13]) );
  DFFR_X1 \Q_reg[12]  ( .D(D[12]), .CK(net18798), .RN(RST), .Q(Q[12]) );
  DFFR_X1 \Q_reg[11]  ( .D(D[11]), .CK(net18798), .RN(RST), .Q(Q[11]) );
  DFFR_X1 \Q_reg[10]  ( .D(D[10]), .CK(net18798), .RN(RST), .Q(Q[10]) );
  DFFR_X1 \Q_reg[9]  ( .D(D[9]), .CK(net18798), .RN(RST), .Q(Q[9]) );
  DFFR_X1 \Q_reg[8]  ( .D(D[8]), .CK(net18798), .RN(RST), .Q(Q[8]) );
  DFFR_X1 \Q_reg[7]  ( .D(D[7]), .CK(net18798), .RN(RST), .Q(Q[7]) );
  DFFR_X1 \Q_reg[6]  ( .D(D[6]), .CK(net18798), .RN(RST), .Q(Q[6]) );
  DFFR_X1 \Q_reg[5]  ( .D(D[5]), .CK(net18798), .RN(RST), .Q(Q[5]) );
  DFFR_X1 \Q_reg[4]  ( .D(D[4]), .CK(net18798), .RN(RST), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(D[3]), .CK(net18798), .RN(RST), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(D[2]), .CK(net18798), .RN(RST), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(D[1]), .CK(net18798), .RN(RST), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(D[0]), .CK(net18798), .RN(RST), .Q(Q[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_reg_N32_4 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18782, net18784, net18786, net18787, net18790, net18793;
  assign net18782 = EN;
  assign net18784 = CLK;
  assign ENCLK = net18786;
  assign net18793 = TE;

  DLL_X1 latch ( .D(net18787), .GN(net18784), .Q(net18790) );
  AND2_X1 main_gate ( .A1(net18790), .A2(net18784), .ZN(net18786) );
  OR2_X1 test_or ( .A1(net18782), .A2(net18793), .ZN(net18787) );
endmodule


module reg_N32_4 ( D, Q, EN, CLK, RST );
  input [31:0] D;
  output [31:0] Q;
  input EN, CLK, RST;
  wire   net18798;

  SNPS_CLOCK_GATE_HIGH_reg_N32_4 clk_gate_Q_reg ( .CLK(CLK), .EN(EN), .ENCLK(
        net18798), .TE(1'b0) );
  DFFR_X1 \Q_reg[31]  ( .D(D[31]), .CK(net18798), .RN(RST), .Q(Q[31]) );
  DFFR_X1 \Q_reg[30]  ( .D(D[30]), .CK(net18798), .RN(RST), .Q(Q[30]) );
  DFFR_X1 \Q_reg[29]  ( .D(D[29]), .CK(net18798), .RN(RST), .Q(Q[29]) );
  DFFR_X1 \Q_reg[28]  ( .D(D[28]), .CK(net18798), .RN(RST), .Q(Q[28]) );
  DFFR_X1 \Q_reg[27]  ( .D(D[27]), .CK(net18798), .RN(RST), .Q(Q[27]) );
  DFFR_X1 \Q_reg[26]  ( .D(D[26]), .CK(net18798), .RN(RST), .Q(Q[26]) );
  DFFR_X1 \Q_reg[25]  ( .D(D[25]), .CK(net18798), .RN(RST), .Q(Q[25]) );
  DFFR_X1 \Q_reg[24]  ( .D(D[24]), .CK(net18798), .RN(RST), .Q(Q[24]) );
  DFFR_X1 \Q_reg[23]  ( .D(D[23]), .CK(net18798), .RN(RST), .Q(Q[23]) );
  DFFR_X1 \Q_reg[22]  ( .D(D[22]), .CK(net18798), .RN(RST), .Q(Q[22]) );
  DFFR_X1 \Q_reg[21]  ( .D(D[21]), .CK(net18798), .RN(RST), .Q(Q[21]) );
  DFFR_X1 \Q_reg[20]  ( .D(D[20]), .CK(net18798), .RN(RST), .Q(Q[20]) );
  DFFR_X1 \Q_reg[19]  ( .D(D[19]), .CK(net18798), .RN(RST), .Q(Q[19]) );
  DFFR_X1 \Q_reg[18]  ( .D(D[18]), .CK(net18798), .RN(RST), .Q(Q[18]) );
  DFFR_X1 \Q_reg[17]  ( .D(D[17]), .CK(net18798), .RN(RST), .Q(Q[17]) );
  DFFR_X1 \Q_reg[16]  ( .D(D[16]), .CK(net18798), .RN(RST), .Q(Q[16]) );
  DFFR_X1 \Q_reg[15]  ( .D(D[15]), .CK(net18798), .RN(RST), .Q(Q[15]) );
  DFFR_X1 \Q_reg[14]  ( .D(D[14]), .CK(net18798), .RN(RST), .Q(Q[14]) );
  DFFR_X1 \Q_reg[13]  ( .D(D[13]), .CK(net18798), .RN(RST), .Q(Q[13]) );
  DFFR_X1 \Q_reg[12]  ( .D(D[12]), .CK(net18798), .RN(RST), .Q(Q[12]) );
  DFFR_X1 \Q_reg[11]  ( .D(D[11]), .CK(net18798), .RN(RST), .Q(Q[11]) );
  DFFR_X1 \Q_reg[10]  ( .D(D[10]), .CK(net18798), .RN(RST), .Q(Q[10]) );
  DFFR_X1 \Q_reg[9]  ( .D(D[9]), .CK(net18798), .RN(RST), .Q(Q[9]) );
  DFFR_X1 \Q_reg[8]  ( .D(D[8]), .CK(net18798), .RN(RST), .Q(Q[8]) );
  DFFR_X1 \Q_reg[7]  ( .D(D[7]), .CK(net18798), .RN(RST), .Q(Q[7]) );
  DFFR_X1 \Q_reg[6]  ( .D(D[6]), .CK(net18798), .RN(RST), .Q(Q[6]) );
  DFFR_X1 \Q_reg[5]  ( .D(D[5]), .CK(net18798), .RN(RST), .Q(Q[5]) );
  DFFR_X1 \Q_reg[4]  ( .D(D[4]), .CK(net18798), .RN(RST), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(D[3]), .CK(net18798), .RN(RST), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(D[2]), .CK(net18798), .RN(RST), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(D[1]), .CK(net18798), .RN(RST), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(D[0]), .CK(net18798), .RN(RST), .Q(Q[0]) );
endmodule


module SNPS_CLOCK_GATE_HIGH_reg_N5_2 ( CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18764, net18766, net18768, net18769, net18772, net18775;
  assign net18764 = EN;
  assign net18766 = CLK;
  assign ENCLK = net18768;
  assign net18775 = TE;

  DLL_X1 latch ( .D(net18769), .GN(net18766), .Q(net18772) );
  AND2_X1 main_gate ( .A1(net18772), .A2(net18766), .ZN(net18768) );
  OR2_X1 test_or ( .A1(net18764), .A2(net18775), .ZN(net18769) );
endmodule


module reg_N5_2 ( D, Q, EN, CLK, RST );
  input [4:0] D;
  output [4:0] Q;
  input EN, CLK, RST;
  wire   net18780;

  SNPS_CLOCK_GATE_HIGH_reg_N5_2 clk_gate_Q_reg ( .CLK(CLK), .EN(EN), .ENCLK(
        net18780), .TE(1'b0) );
  DFFR_X1 \Q_reg[4]  ( .D(D[4]), .CK(net18780), .RN(RST), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(D[3]), .CK(net18780), .RN(RST), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(D[2]), .CK(net18780), .RN(RST), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(D[1]), .CK(net18780), .RN(RST), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(D[0]), .CK(net18780), .RN(RST), .Q(Q[0]) );
endmodule


module MUX_8to1_N32_2 ( IN0, IN1, IN2, IN3, IN4, IN5, IN6, IN7, SEL, Y );
  input [31:0] IN0;
  input [31:0] IN1;
  input [31:0] IN2;
  input [31:0] IN3;
  input [31:0] IN4;
  input [31:0] IN5;
  input [31:0] IN6;
  input [31:0] IN7;
  input [2:0] SEL;
  output [31:0] Y;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32;

  AND2_X1 U1 ( .A1(IN4[3]), .A2(n1), .ZN(Y[3]) );
  AND2_X1 U2 ( .A1(IN4[2]), .A2(n1), .ZN(Y[2]) );
  AND2_X1 U3 ( .A1(IN0[8]), .A2(n1), .ZN(Y[7]) );
  AOI21_X1 U4 ( .B1(SEL[1]), .B2(n12), .A(n31), .ZN(n11) );
  AND2_X1 U5 ( .A1(IN4[4]), .A2(n1), .ZN(Y[4]) );
  AND2_X1 U6 ( .A1(IN4[0]), .A2(n1), .ZN(Y[0]) );
  AND2_X1 U7 ( .A1(IN4[6]), .A2(n1), .ZN(Y[6]) );
  AND2_X1 U8 ( .A1(IN4[5]), .A2(n1), .ZN(Y[5]) );
  AND2_X1 U9 ( .A1(IN4[1]), .A2(n1), .ZN(Y[1]) );
  OR2_X1 U10 ( .A1(n12), .A2(n2), .ZN(n1) );
  NAND3_X1 U11 ( .A1(n2), .A2(IN0[8]), .A3(n12), .ZN(n13) );
  INV_X1 U12 ( .A(SEL[2]), .ZN(n12) );
  OAI21_X2 U13 ( .B1(SEL[0]), .B2(n14), .A(n13), .ZN(n30) );
  NOR3_X4 U14 ( .A1(SEL[1]), .A2(SEL[0]), .A3(n12), .ZN(n31) );
  NOR2_X1 U15 ( .A1(SEL[1]), .A2(SEL[0]), .ZN(n2) );
  INV_X1 U16 ( .A(IN4[8]), .ZN(n3) );
  OAI21_X1 U17 ( .B1(n11), .B2(n3), .A(n13), .ZN(Y[8]) );
  INV_X1 U18 ( .A(IN4[9]), .ZN(n4) );
  OAI21_X1 U19 ( .B1(n11), .B2(n4), .A(n13), .ZN(Y[9]) );
  INV_X1 U20 ( .A(IN4[10]), .ZN(n5) );
  OAI21_X1 U21 ( .B1(n11), .B2(n5), .A(n13), .ZN(Y[10]) );
  INV_X1 U22 ( .A(IN4[11]), .ZN(n6) );
  OAI21_X1 U23 ( .B1(n11), .B2(n6), .A(n13), .ZN(Y[11]) );
  INV_X1 U24 ( .A(IN4[12]), .ZN(n7) );
  OAI21_X1 U25 ( .B1(n11), .B2(n7), .A(n13), .ZN(Y[12]) );
  INV_X1 U26 ( .A(IN4[13]), .ZN(n8) );
  OAI21_X1 U27 ( .B1(n11), .B2(n8), .A(n13), .ZN(Y[13]) );
  INV_X1 U28 ( .A(IN4[14]), .ZN(n9) );
  OAI21_X1 U29 ( .B1(n11), .B2(n9), .A(n13), .ZN(Y[14]) );
  INV_X1 U30 ( .A(IN2[16]), .ZN(n10) );
  OAI21_X1 U31 ( .B1(n11), .B2(n10), .A(n13), .ZN(Y[15]) );
  NAND3_X1 U32 ( .A1(SEL[1]), .A2(IN2[16]), .A3(n12), .ZN(n14) );
  AOI21_X1 U33 ( .B1(n31), .B2(IN4[16]), .A(n30), .ZN(n15) );
  INV_X1 U34 ( .A(n15), .ZN(Y[16]) );
  AOI21_X1 U35 ( .B1(n31), .B2(IN4[17]), .A(n30), .ZN(n16) );
  INV_X1 U36 ( .A(n16), .ZN(Y[17]) );
  AOI21_X1 U37 ( .B1(n31), .B2(IN4[18]), .A(n30), .ZN(n17) );
  INV_X1 U38 ( .A(n17), .ZN(Y[18]) );
  AOI21_X1 U39 ( .B1(n31), .B2(IN4[19]), .A(n30), .ZN(n18) );
  INV_X1 U40 ( .A(n18), .ZN(Y[19]) );
  AOI21_X1 U41 ( .B1(n31), .B2(IN4[20]), .A(n30), .ZN(n19) );
  INV_X1 U42 ( .A(n19), .ZN(Y[20]) );
  AOI21_X1 U43 ( .B1(n31), .B2(IN4[21]), .A(n30), .ZN(n20) );
  INV_X1 U44 ( .A(n20), .ZN(Y[21]) );
  AOI21_X1 U45 ( .B1(n31), .B2(IN4[22]), .A(n30), .ZN(n21) );
  INV_X1 U46 ( .A(n21), .ZN(Y[22]) );
  AOI21_X1 U47 ( .B1(n31), .B2(IN4[23]), .A(n30), .ZN(n22) );
  INV_X1 U48 ( .A(n22), .ZN(Y[23]) );
  AOI21_X1 U49 ( .B1(n31), .B2(IN4[24]), .A(n30), .ZN(n23) );
  INV_X1 U50 ( .A(n23), .ZN(Y[24]) );
  AOI21_X1 U51 ( .B1(n31), .B2(IN4[25]), .A(n30), .ZN(n24) );
  INV_X1 U52 ( .A(n24), .ZN(Y[25]) );
  AOI21_X1 U53 ( .B1(n31), .B2(IN4[26]), .A(n30), .ZN(n25) );
  INV_X1 U54 ( .A(n25), .ZN(Y[26]) );
  AOI21_X1 U55 ( .B1(n31), .B2(IN4[27]), .A(n30), .ZN(n26) );
  INV_X1 U56 ( .A(n26), .ZN(Y[27]) );
  AOI21_X1 U57 ( .B1(n31), .B2(IN4[28]), .A(n30), .ZN(n27) );
  INV_X1 U58 ( .A(n27), .ZN(Y[28]) );
  AOI21_X1 U59 ( .B1(n31), .B2(IN4[29]), .A(n30), .ZN(n28) );
  INV_X1 U60 ( .A(n28), .ZN(Y[29]) );
  AOI21_X1 U61 ( .B1(n31), .B2(IN4[30]), .A(n30), .ZN(n29) );
  INV_X1 U62 ( .A(n29), .ZN(Y[30]) );
  AOI21_X1 U63 ( .B1(n31), .B2(IN4[31]), .A(n30), .ZN(n32) );
  INV_X1 U64 ( .A(n32), .ZN(Y[31]) );
endmodule


module reg_N32_3 ( D, Q, EN, CLK, RST );
  input [31:0] D;
  output [31:0] Q;
  input EN, CLK, RST;


  DFFR_X1 \Q_reg[31]  ( .D(D[31]), .CK(CLK), .RN(RST), .Q(Q[31]) );
  DFFR_X1 \Q_reg[30]  ( .D(D[30]), .CK(CLK), .RN(RST), .Q(Q[30]) );
  DFFR_X1 \Q_reg[29]  ( .D(D[29]), .CK(CLK), .RN(RST), .Q(Q[29]) );
  DFFR_X1 \Q_reg[28]  ( .D(D[28]), .CK(CLK), .RN(RST), .Q(Q[28]) );
  DFFR_X1 \Q_reg[27]  ( .D(D[27]), .CK(CLK), .RN(RST), .Q(Q[27]) );
  DFFR_X1 \Q_reg[26]  ( .D(D[26]), .CK(CLK), .RN(RST), .Q(Q[26]) );
  DFFR_X1 \Q_reg[25]  ( .D(D[25]), .CK(CLK), .RN(RST), .Q(Q[25]) );
  DFFR_X1 \Q_reg[24]  ( .D(D[24]), .CK(CLK), .RN(RST), .Q(Q[24]) );
  DFFR_X1 \Q_reg[23]  ( .D(D[23]), .CK(CLK), .RN(RST), .Q(Q[23]) );
  DFFR_X1 \Q_reg[22]  ( .D(D[22]), .CK(CLK), .RN(RST), .Q(Q[22]) );
  DFFR_X1 \Q_reg[21]  ( .D(D[21]), .CK(CLK), .RN(RST), .Q(Q[21]) );
  DFFR_X1 \Q_reg[20]  ( .D(D[20]), .CK(CLK), .RN(RST), .Q(Q[20]) );
  DFFR_X1 \Q_reg[19]  ( .D(D[19]), .CK(CLK), .RN(RST), .Q(Q[19]) );
  DFFR_X1 \Q_reg[18]  ( .D(D[18]), .CK(CLK), .RN(RST), .Q(Q[18]) );
  DFFR_X1 \Q_reg[17]  ( .D(D[17]), .CK(CLK), .RN(RST), .Q(Q[17]) );
  DFFR_X1 \Q_reg[16]  ( .D(D[16]), .CK(CLK), .RN(RST), .Q(Q[16]) );
  DFFR_X1 \Q_reg[15]  ( .D(D[15]), .CK(CLK), .RN(RST), .Q(Q[15]) );
  DFFR_X1 \Q_reg[14]  ( .D(D[14]), .CK(CLK), .RN(RST), .Q(Q[14]) );
  DFFR_X1 \Q_reg[13]  ( .D(D[13]), .CK(CLK), .RN(RST), .Q(Q[13]) );
  DFFR_X1 \Q_reg[12]  ( .D(D[12]), .CK(CLK), .RN(RST), .Q(Q[12]) );
  DFFR_X1 \Q_reg[11]  ( .D(D[11]), .CK(CLK), .RN(RST), .Q(Q[11]) );
  DFFR_X1 \Q_reg[10]  ( .D(D[10]), .CK(CLK), .RN(RST), .Q(Q[10]) );
  DFFR_X1 \Q_reg[9]  ( .D(D[9]), .CK(CLK), .RN(RST), .Q(Q[9]) );
  DFFR_X1 \Q_reg[8]  ( .D(D[8]), .CK(CLK), .RN(RST), .Q(Q[8]) );
  DFFR_X1 \Q_reg[7]  ( .D(D[7]), .CK(CLK), .RN(RST), .Q(Q[7]) );
  DFFR_X1 \Q_reg[6]  ( .D(D[6]), .CK(CLK), .RN(RST), .Q(Q[6]) );
  DFFR_X1 \Q_reg[5]  ( .D(D[5]), .CK(CLK), .RN(RST), .Q(Q[5]) );
  DFFR_X1 \Q_reg[4]  ( .D(D[4]), .CK(CLK), .RN(RST), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(D[3]), .CK(CLK), .RN(RST), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(D[2]), .CK(CLK), .RN(RST), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(D[1]), .CK(CLK), .RN(RST), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(D[0]), .CK(CLK), .RN(RST), .Q(Q[0]) );
endmodule


module reg_N32_2 ( D, Q, EN, CLK, RST );
  input [31:0] D;
  output [31:0] Q;
  input EN, CLK, RST;


  DFFR_X1 \Q_reg[31]  ( .D(D[31]), .CK(CLK), .RN(RST), .Q(Q[31]) );
  DFFR_X1 \Q_reg[30]  ( .D(D[30]), .CK(CLK), .RN(RST), .Q(Q[30]) );
  DFFR_X1 \Q_reg[29]  ( .D(D[29]), .CK(CLK), .RN(RST), .Q(Q[29]) );
  DFFR_X1 \Q_reg[28]  ( .D(D[28]), .CK(CLK), .RN(RST), .Q(Q[28]) );
  DFFR_X1 \Q_reg[27]  ( .D(D[27]), .CK(CLK), .RN(RST), .Q(Q[27]) );
  DFFR_X1 \Q_reg[26]  ( .D(D[26]), .CK(CLK), .RN(RST), .Q(Q[26]) );
  DFFR_X1 \Q_reg[25]  ( .D(D[25]), .CK(CLK), .RN(RST), .Q(Q[25]) );
  DFFR_X1 \Q_reg[24]  ( .D(D[24]), .CK(CLK), .RN(RST), .Q(Q[24]) );
  DFFR_X1 \Q_reg[23]  ( .D(D[23]), .CK(CLK), .RN(RST), .Q(Q[23]) );
  DFFR_X1 \Q_reg[22]  ( .D(D[22]), .CK(CLK), .RN(RST), .Q(Q[22]) );
  DFFR_X1 \Q_reg[21]  ( .D(D[21]), .CK(CLK), .RN(RST), .Q(Q[21]) );
  DFFR_X1 \Q_reg[20]  ( .D(D[20]), .CK(CLK), .RN(RST), .Q(Q[20]) );
  DFFR_X1 \Q_reg[19]  ( .D(D[19]), .CK(CLK), .RN(RST), .Q(Q[19]) );
  DFFR_X1 \Q_reg[18]  ( .D(D[18]), .CK(CLK), .RN(RST), .Q(Q[18]) );
  DFFR_X1 \Q_reg[17]  ( .D(D[17]), .CK(CLK), .RN(RST), .Q(Q[17]) );
  DFFR_X1 \Q_reg[16]  ( .D(D[16]), .CK(CLK), .RN(RST), .Q(Q[16]) );
  DFFR_X1 \Q_reg[15]  ( .D(D[15]), .CK(CLK), .RN(RST), .Q(Q[15]) );
  DFFR_X1 \Q_reg[14]  ( .D(D[14]), .CK(CLK), .RN(RST), .Q(Q[14]) );
  DFFR_X1 \Q_reg[13]  ( .D(D[13]), .CK(CLK), .RN(RST), .Q(Q[13]) );
  DFFR_X1 \Q_reg[12]  ( .D(D[12]), .CK(CLK), .RN(RST), .Q(Q[12]) );
  DFFR_X1 \Q_reg[11]  ( .D(D[11]), .CK(CLK), .RN(RST), .Q(Q[11]) );
  DFFR_X1 \Q_reg[10]  ( .D(D[10]), .CK(CLK), .RN(RST), .Q(Q[10]) );
  DFFR_X1 \Q_reg[9]  ( .D(D[9]), .CK(CLK), .RN(RST), .Q(Q[9]) );
  DFFR_X1 \Q_reg[8]  ( .D(D[8]), .CK(CLK), .RN(RST), .Q(Q[8]) );
  DFFR_X1 \Q_reg[7]  ( .D(D[7]), .CK(CLK), .RN(RST), .Q(Q[7]) );
  DFFR_X1 \Q_reg[6]  ( .D(D[6]), .CK(CLK), .RN(RST), .Q(Q[6]) );
  DFFR_X1 \Q_reg[5]  ( .D(D[5]), .CK(CLK), .RN(RST), .Q(Q[5]) );
  DFFR_X1 \Q_reg[4]  ( .D(D[4]), .CK(CLK), .RN(RST), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(D[3]), .CK(CLK), .RN(RST), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(D[2]), .CK(CLK), .RN(RST), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(D[1]), .CK(CLK), .RN(RST), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(D[0]), .CK(CLK), .RN(RST), .Q(Q[0]) );
endmodule


module reg_N32_1 ( D, Q, EN, CLK, RST );
  input [31:0] D;
  output [31:0] Q;
  input EN, CLK, RST;


  DFFR_X1 \Q_reg[31]  ( .D(D[31]), .CK(CLK), .RN(RST), .Q(Q[31]) );
  DFFR_X1 \Q_reg[30]  ( .D(D[30]), .CK(CLK), .RN(RST), .Q(Q[30]) );
  DFFR_X1 \Q_reg[29]  ( .D(D[29]), .CK(CLK), .RN(RST), .Q(Q[29]) );
  DFFR_X1 \Q_reg[28]  ( .D(D[28]), .CK(CLK), .RN(RST), .Q(Q[28]) );
  DFFR_X1 \Q_reg[27]  ( .D(D[27]), .CK(CLK), .RN(RST), .Q(Q[27]) );
  DFFR_X1 \Q_reg[26]  ( .D(D[26]), .CK(CLK), .RN(RST), .Q(Q[26]) );
  DFFR_X1 \Q_reg[25]  ( .D(D[25]), .CK(CLK), .RN(RST), .Q(Q[25]) );
  DFFR_X1 \Q_reg[24]  ( .D(D[24]), .CK(CLK), .RN(RST), .Q(Q[24]) );
  DFFR_X1 \Q_reg[23]  ( .D(D[23]), .CK(CLK), .RN(RST), .Q(Q[23]) );
  DFFR_X1 \Q_reg[22]  ( .D(D[22]), .CK(CLK), .RN(RST), .Q(Q[22]) );
  DFFR_X1 \Q_reg[21]  ( .D(D[21]), .CK(CLK), .RN(RST), .Q(Q[21]) );
  DFFR_X1 \Q_reg[20]  ( .D(D[20]), .CK(CLK), .RN(RST), .Q(Q[20]) );
  DFFR_X1 \Q_reg[19]  ( .D(D[19]), .CK(CLK), .RN(RST), .Q(Q[19]) );
  DFFR_X1 \Q_reg[18]  ( .D(D[18]), .CK(CLK), .RN(RST), .Q(Q[18]) );
  DFFR_X1 \Q_reg[17]  ( .D(D[17]), .CK(CLK), .RN(RST), .Q(Q[17]) );
  DFFR_X1 \Q_reg[16]  ( .D(D[16]), .CK(CLK), .RN(RST), .Q(Q[16]) );
  DFFR_X1 \Q_reg[15]  ( .D(D[15]), .CK(CLK), .RN(RST), .Q(Q[15]) );
  DFFR_X1 \Q_reg[14]  ( .D(D[14]), .CK(CLK), .RN(RST), .Q(Q[14]) );
  DFFR_X1 \Q_reg[13]  ( .D(D[13]), .CK(CLK), .RN(RST), .Q(Q[13]) );
  DFFR_X1 \Q_reg[12]  ( .D(D[12]), .CK(CLK), .RN(RST), .Q(Q[12]) );
  DFFR_X1 \Q_reg[11]  ( .D(D[11]), .CK(CLK), .RN(RST), .Q(Q[11]) );
  DFFR_X1 \Q_reg[10]  ( .D(D[10]), .CK(CLK), .RN(RST), .Q(Q[10]) );
  DFFR_X1 \Q_reg[9]  ( .D(D[9]), .CK(CLK), .RN(RST), .Q(Q[9]) );
  DFFR_X1 \Q_reg[8]  ( .D(D[8]), .CK(CLK), .RN(RST), .Q(Q[8]) );
  DFFR_X1 \Q_reg[7]  ( .D(D[7]), .CK(CLK), .RN(RST), .Q(Q[7]) );
  DFFR_X1 \Q_reg[6]  ( .D(D[6]), .CK(CLK), .RN(RST), .Q(Q[6]) );
  DFFR_X1 \Q_reg[5]  ( .D(D[5]), .CK(CLK), .RN(RST), .Q(Q[5]) );
  DFFR_X1 \Q_reg[4]  ( .D(D[4]), .CK(CLK), .RN(RST), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(D[3]), .CK(CLK), .RN(RST), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(D[2]), .CK(CLK), .RN(RST), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(D[1]), .CK(CLK), .RN(RST), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(D[0]), .CK(CLK), .RN(RST), .Q(Q[0]) );
endmodule


module reg_N5_1 ( D, Q, EN, CLK, RST );
  input [4:0] D;
  output [4:0] Q;
  input EN, CLK, RST;


  DFFR_X1 \Q_reg[4]  ( .D(D[4]), .CK(CLK), .RN(RST), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(D[3]), .CK(CLK), .RN(RST), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(D[2]), .CK(CLK), .RN(RST), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(D[1]), .CK(CLK), .RN(RST), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(D[0]), .CK(CLK), .RN(RST), .Q(Q[0]) );
endmodule


module MUX_4to1_N32 ( IN0, IN1, IN2, IN3, SEL, Y );
  input [31:0] IN0;
  input [31:0] IN1;
  input [31:0] IN2;
  input [31:0] IN3;
  input [1:0] SEL;
  output [31:0] Y;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38;

  INV_X2 U1 ( .A(n9), .ZN(Y[14]) );
  INV_X2 U2 ( .A(n4), .ZN(Y[0]) );
  INV_X2 U3 ( .A(n19), .ZN(Y[23]) );
  INV_X2 U4 ( .A(n26), .ZN(Y[2]) );
  INV_X2 U5 ( .A(n28), .ZN(Y[31]) );
  INV_X2 U6 ( .A(n34), .ZN(Y[8]) );
  INV_X2 U7 ( .A(n31), .ZN(Y[5]) );
  INV_X2 U8 ( .A(n33), .ZN(Y[7]) );
  INV_X2 U9 ( .A(n32), .ZN(Y[6]) );
  INV_X2 U10 ( .A(n27), .ZN(Y[30]) );
  INV_X2 U11 ( .A(n5), .ZN(Y[10]) );
  INV_X2 U12 ( .A(n30), .ZN(Y[4]) );
  INV_X2 U13 ( .A(n38), .ZN(Y[9]) );
  INV_X2 U14 ( .A(n23), .ZN(Y[27]) );
  INV_X2 U15 ( .A(n15), .ZN(Y[1]) );
  INV_X2 U16 ( .A(n18), .ZN(Y[22]) );
  INV_X2 U17 ( .A(n8), .ZN(Y[13]) );
  INV_X2 U18 ( .A(n16), .ZN(Y[20]) );
  INV_X2 U19 ( .A(n29), .ZN(Y[3]) );
  INV_X2 U20 ( .A(n17), .ZN(Y[21]) );
  INV_X2 U21 ( .A(n14), .ZN(Y[19]) );
  INV_X2 U22 ( .A(n22), .ZN(Y[26]) );
  INV_X2 U23 ( .A(n20), .ZN(Y[24]) );
  INV_X2 U24 ( .A(n11), .ZN(Y[16]) );
  INV_X2 U25 ( .A(n13), .ZN(Y[18]) );
  INV_X2 U26 ( .A(n25), .ZN(Y[29]) );
  INV_X2 U27 ( .A(n6), .ZN(Y[11]) );
  INV_X2 U28 ( .A(n24), .ZN(Y[28]) );
  INV_X2 U29 ( .A(n10), .ZN(Y[15]) );
  INV_X2 U30 ( .A(n12), .ZN(Y[17]) );
  INV_X2 U31 ( .A(n21), .ZN(Y[25]) );
  INV_X2 U32 ( .A(n7), .ZN(Y[12]) );
  NOR2_X1 U33 ( .A1(SEL[1]), .A2(SEL[0]), .ZN(n35) );
  BUF_X1 U34 ( .A(n36), .Z(n2) );
  BUF_X1 U35 ( .A(n35), .Z(n1) );
  NOR2_X1 U36 ( .A1(SEL[0]), .A2(n3), .ZN(n36) );
  AND2_X2 U37 ( .A1(n3), .A2(SEL[0]), .ZN(n37) );
  INV_X1 U38 ( .A(SEL[1]), .ZN(n3) );
  AOI222_X1 U39 ( .A1(n37), .A2(IN1[0]), .B1(n2), .B2(IN2[0]), .C1(n1), .C2(
        IN0[0]), .ZN(n4) );
  AOI222_X1 U40 ( .A1(n37), .A2(IN1[10]), .B1(n2), .B2(IN2[10]), .C1(n1), .C2(
        IN0[10]), .ZN(n5) );
  AOI222_X1 U41 ( .A1(n37), .A2(IN1[11]), .B1(n36), .B2(IN2[11]), .C1(n35), 
        .C2(IN0[11]), .ZN(n6) );
  AOI222_X1 U42 ( .A1(n37), .A2(IN1[12]), .B1(n36), .B2(IN2[12]), .C1(n35), 
        .C2(IN0[12]), .ZN(n7) );
  AOI222_X1 U43 ( .A1(n37), .A2(IN1[13]), .B1(n2), .B2(IN2[13]), .C1(n1), .C2(
        IN0[13]), .ZN(n8) );
  AOI222_X1 U44 ( .A1(n37), .A2(IN1[14]), .B1(n2), .B2(IN2[14]), .C1(n1), .C2(
        IN0[14]), .ZN(n9) );
  AOI222_X1 U45 ( .A1(n37), .A2(IN1[15]), .B1(n36), .B2(IN2[15]), .C1(n35), 
        .C2(IN0[15]), .ZN(n10) );
  AOI222_X1 U46 ( .A1(n37), .A2(IN1[16]), .B1(n36), .B2(IN2[16]), .C1(n35), 
        .C2(IN0[16]), .ZN(n11) );
  AOI222_X1 U47 ( .A1(n37), .A2(IN1[17]), .B1(n36), .B2(IN2[17]), .C1(n35), 
        .C2(IN0[17]), .ZN(n12) );
  AOI222_X1 U48 ( .A1(n37), .A2(IN1[18]), .B1(n36), .B2(IN2[18]), .C1(n35), 
        .C2(IN0[18]), .ZN(n13) );
  AOI222_X1 U49 ( .A1(n37), .A2(IN1[19]), .B1(n2), .B2(IN2[19]), .C1(n1), .C2(
        IN0[19]), .ZN(n14) );
  AOI222_X1 U50 ( .A1(n37), .A2(IN1[1]), .B1(n2), .B2(IN2[1]), .C1(n35), .C2(
        IN0[1]), .ZN(n15) );
  AOI222_X1 U51 ( .A1(n37), .A2(IN1[20]), .B1(n2), .B2(IN2[20]), .C1(n35), 
        .C2(IN0[20]), .ZN(n16) );
  AOI222_X1 U52 ( .A1(n37), .A2(IN1[21]), .B1(n2), .B2(IN2[21]), .C1(n1), .C2(
        IN0[21]), .ZN(n17) );
  AOI222_X1 U53 ( .A1(n37), .A2(IN1[22]), .B1(n2), .B2(IN2[22]), .C1(n35), 
        .C2(IN0[22]), .ZN(n18) );
  AOI222_X1 U54 ( .A1(n37), .A2(IN1[23]), .B1(n2), .B2(IN2[23]), .C1(n1), .C2(
        IN0[23]), .ZN(n19) );
  AOI222_X1 U55 ( .A1(n37), .A2(IN1[24]), .B1(n36), .B2(IN2[24]), .C1(n1), 
        .C2(IN0[24]), .ZN(n20) );
  AOI222_X1 U56 ( .A1(n37), .A2(IN1[25]), .B1(n36), .B2(IN2[25]), .C1(n1), 
        .C2(IN0[25]), .ZN(n21) );
  AOI222_X1 U57 ( .A1(n37), .A2(IN1[26]), .B1(n2), .B2(IN2[26]), .C1(n35), 
        .C2(IN0[26]), .ZN(n22) );
  AOI222_X1 U58 ( .A1(n37), .A2(IN1[27]), .B1(n2), .B2(IN2[27]), .C1(n35), 
        .C2(IN0[27]), .ZN(n23) );
  AOI222_X1 U59 ( .A1(n37), .A2(IN1[28]), .B1(n36), .B2(IN2[28]), .C1(n1), 
        .C2(IN0[28]), .ZN(n24) );
  AOI222_X1 U60 ( .A1(n37), .A2(IN1[29]), .B1(n36), .B2(IN2[29]), .C1(n1), 
        .C2(IN0[29]), .ZN(n25) );
  AOI222_X1 U61 ( .A1(n37), .A2(IN1[2]), .B1(n2), .B2(IN2[2]), .C1(n1), .C2(
        IN0[2]), .ZN(n26) );
  AOI222_X1 U62 ( .A1(n37), .A2(IN1[30]), .B1(n2), .B2(IN2[30]), .C1(n1), .C2(
        IN0[30]), .ZN(n27) );
  AOI222_X1 U63 ( .A1(n37), .A2(IN1[31]), .B1(n2), .B2(IN2[31]), .C1(n1), .C2(
        IN0[31]), .ZN(n28) );
  AOI222_X1 U64 ( .A1(n37), .A2(IN1[3]), .B1(n2), .B2(IN2[3]), .C1(n1), .C2(
        IN0[3]), .ZN(n29) );
  AOI222_X1 U65 ( .A1(n37), .A2(IN1[4]), .B1(n2), .B2(IN2[4]), .C1(n1), .C2(
        IN0[4]), .ZN(n30) );
  AOI222_X1 U66 ( .A1(n37), .A2(IN1[5]), .B1(n2), .B2(IN2[5]), .C1(n1), .C2(
        IN0[5]), .ZN(n31) );
  AOI222_X1 U67 ( .A1(n37), .A2(IN1[6]), .B1(n2), .B2(IN2[6]), .C1(n1), .C2(
        IN0[6]), .ZN(n32) );
  AOI222_X1 U68 ( .A1(n37), .A2(IN1[7]), .B1(n2), .B2(IN2[7]), .C1(n1), .C2(
        IN0[7]), .ZN(n33) );
  AOI222_X1 U69 ( .A1(n37), .A2(IN1[8]), .B1(n2), .B2(IN2[8]), .C1(n1), .C2(
        IN0[8]), .ZN(n34) );
  AOI222_X1 U70 ( .A1(n37), .A2(IN1[9]), .B1(n2), .B2(IN2[9]), .C1(n1), .C2(
        IN0[9]), .ZN(n38) );
endmodule


module datapath_BPU_TAG_FIELD_SIZE8_BPU_SET_FIELD_SIZE3_BPU_LINES_PER_SET4 ( 
        IRAM_OUT, DRAM_ADDR, DRAM_IN, DRAM_OUT, .control_from_CU({
        \control_from_CU[ID][MUX_BRANCH_SEL] , 
        \control_from_CU[ID][MUX_IMM_EXT_SEL] , 
        \control_from_CU[ID][MUX_RF_WR_ADDR_SEL][1] , 
        \control_from_CU[ID][MUX_RF_WR_ADDR_SEL][0] , 
        \control_from_CU[ID][BRANCH_COND][1] , 
        \control_from_CU[ID][BRANCH_COND][0] , \control_from_CU[EXE][MULT_EN] , 
        \control_from_CU[EXE][MUX_MULT_SEL] , 
        \control_from_CU[EXE][MUX_ALU_IN2_SEL] , 
        \control_from_CU[EXE][ALU_OP][4] , \control_from_CU[EXE][ALU_OP][3] , 
        \control_from_CU[EXE][ALU_OP][2] , \control_from_CU[EXE][ALU_OP][1] , 
        \control_from_CU[EXE][ALU_OP][0] , 
        \control_from_CU[MEM][DRAM_WR_EN][1] , 
        \control_from_CU[MEM][DRAM_WR_EN][0] , 
        \control_from_CU[MEM][MUX_DRAM_OUT_EXT_SEL][2] , 
        \control_from_CU[MEM][MUX_DRAM_OUT_EXT_SEL][1] , 
        \control_from_CU[MEM][MUX_DRAM_OUT_EXT_SEL][0] , 
        \control_from_CU[WB][MUX_WB_SEL][1] , 
        \control_from_CU[WB][MUX_WB_SEL][0] , \control_from_CU[WB][RF_WR_EN] }
        ), .control_from_FU({\control_from_FU[MUX_RF_OUT1_SEL][2] , 
        \control_from_FU[MUX_RF_OUT1_SEL][1] , 
        \control_from_FU[MUX_RF_OUT1_SEL][0] , 
        \control_from_FU[MUX_RF_OUT2_SEL][2] , 
        \control_from_FU[MUX_RF_OUT2_SEL][1] , 
        \control_from_FU[MUX_RF_OUT2_SEL][0] , 
        \control_from_FU[MUX_DRAM_IN_SEL] }), .control_from_HDU({
        \control_from_HDU[PC_EN] , \control_from_HDU[IF_EN] , 
        \control_from_HDU[ID_EN] , \control_from_HDU[EXE_EN] , 
        \control_from_HDU[MEM_EN] , \control_from_HDU[WB_EN] , 
        \control_from_HDU[ID_BUBBLE] , \control_from_HDU[EXE_BUBBLE] , 
        \control_from_HDU[MEM_BUBBLE] , \control_from_HDU[WB_BUBBLE] }), CLK, 
        RST, \IRAM_ADDR[31] , \IRAM_ADDR[30] , \IRAM_ADDR[29] , 
        \IRAM_ADDR[28] , \IRAM_ADDR[27] , \IRAM_ADDR[26] , \IRAM_ADDR[25] , 
        \IRAM_ADDR[24] , \IRAM_ADDR[23] , \IRAM_ADDR[22] , \IRAM_ADDR[21] , 
        \IRAM_ADDR[20] , \IRAM_ADDR[19] , \IRAM_ADDR[18] , \IRAM_ADDR[17] , 
        \IRAM_ADDR[16] , \IRAM_ADDR[15] , \IRAM_ADDR[14] , \IRAM_ADDR[13] , 
        \IRAM_ADDR[12] , \IRAM_ADDR[11] , \IRAM_ADDR[10] , \IRAM_ADDR[9] , 
        \IRAM_ADDR[8] , \IRAM_ADDR[7] , \IRAM_ADDR[6] , \IRAM_ADDR[5] , 
        \IRAM_ADDR[1] , \IRAM_ADDR[0] , \IRAM_ADDR[3]_BAR , misprediction_BAR, 
        \IRAM_ADDR[2] , \IRAM_ADDR[4]_BAR  );
  input [31:0] IRAM_OUT;
  output [31:0] DRAM_ADDR;
  output [31:0] DRAM_IN;
  input [31:0] DRAM_OUT;
  input \control_from_CU[ID][MUX_BRANCH_SEL] ,
         \control_from_CU[ID][MUX_IMM_EXT_SEL] ,
         \control_from_CU[ID][MUX_RF_WR_ADDR_SEL][1] ,
         \control_from_CU[ID][MUX_RF_WR_ADDR_SEL][0] ,
         \control_from_CU[ID][BRANCH_COND][1] ,
         \control_from_CU[ID][BRANCH_COND][0] ,
         \control_from_CU[EXE][MULT_EN] , \control_from_CU[EXE][MUX_MULT_SEL] ,
         \control_from_CU[EXE][MUX_ALU_IN2_SEL] ,
         \control_from_CU[EXE][ALU_OP][4] , \control_from_CU[EXE][ALU_OP][3] ,
         \control_from_CU[EXE][ALU_OP][2] , \control_from_CU[EXE][ALU_OP][1] ,
         \control_from_CU[EXE][ALU_OP][0] ,
         \control_from_CU[MEM][DRAM_WR_EN][1] ,
         \control_from_CU[MEM][DRAM_WR_EN][0] ,
         \control_from_CU[MEM][MUX_DRAM_OUT_EXT_SEL][2] ,
         \control_from_CU[MEM][MUX_DRAM_OUT_EXT_SEL][1] ,
         \control_from_CU[MEM][MUX_DRAM_OUT_EXT_SEL][0] ,
         \control_from_CU[WB][MUX_WB_SEL][1] ,
         \control_from_CU[WB][MUX_WB_SEL][0] , \control_from_CU[WB][RF_WR_EN] ,
         \control_from_FU[MUX_RF_OUT1_SEL][2] ,
         \control_from_FU[MUX_RF_OUT1_SEL][1] ,
         \control_from_FU[MUX_RF_OUT1_SEL][0] ,
         \control_from_FU[MUX_RF_OUT2_SEL][2] ,
         \control_from_FU[MUX_RF_OUT2_SEL][1] ,
         \control_from_FU[MUX_RF_OUT2_SEL][0] ,
         \control_from_FU[MUX_DRAM_IN_SEL] , \control_from_HDU[PC_EN] ,
         \control_from_HDU[IF_EN] , \control_from_HDU[ID_EN] ,
         \control_from_HDU[EXE_EN] , \control_from_HDU[MEM_EN] ,
         \control_from_HDU[WB_EN] , \control_from_HDU[ID_BUBBLE] ,
         \control_from_HDU[EXE_BUBBLE] , \control_from_HDU[MEM_BUBBLE] ,
         \control_from_HDU[WB_BUBBLE] , CLK, RST;
  output \IRAM_ADDR[31] , \IRAM_ADDR[30] , \IRAM_ADDR[29] , \IRAM_ADDR[28] ,
         \IRAM_ADDR[27] , \IRAM_ADDR[26] , \IRAM_ADDR[25] , \IRAM_ADDR[24] ,
         \IRAM_ADDR[23] , \IRAM_ADDR[22] , \IRAM_ADDR[21] , \IRAM_ADDR[20] ,
         \IRAM_ADDR[19] , \IRAM_ADDR[18] , \IRAM_ADDR[17] , \IRAM_ADDR[16] ,
         \IRAM_ADDR[15] , \IRAM_ADDR[14] , \IRAM_ADDR[13] , \IRAM_ADDR[12] ,
         \IRAM_ADDR[11] , \IRAM_ADDR[10] , \IRAM_ADDR[9] , \IRAM_ADDR[8] ,
         \IRAM_ADDR[7] , \IRAM_ADDR[6] , \IRAM_ADDR[5] , \IRAM_ADDR[1] ,
         \IRAM_ADDR[0] , \IRAM_ADDR[3]_BAR , misprediction_BAR, \IRAM_ADDR[2] ,
         \IRAM_ADDR[4]_BAR ;
  wire   misprediction, branch_is_taken, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n155, n156, n157;
  wire   [31:0] IRAM_ADDR;
  wire   [31:0] PC_IN;
  wire   [31:0] NPC;
  wire   [31:0] actual_addr;
  wire   [31:0] NPC_ID;
  wire   [25:0] IR_out;
  wire   [31:0] RF_OUT1_fw;
  wire   [31:0] ADDER_BRANCH_out;
  wire   [31:0] NPC_BRANCH;
  wire   [31:0] IMM_ID;
  wire   [31:0] RF_OUT1;
  wire   [31:0] ALU_OUT_EXE;
  wire   [31:0] LMD_in;
  wire   [31:0] NPC_MEM;
  wire   [31:0] NPC_EXE;
  wire   [31:0] RF_OUT2;
  wire   [31:0] RF_OUT2_fw;
  wire   [4:0] RF_WR_ADDR_ID;
  wire   [4:0] RF_WR_ADDR_EXE;
  wire   [4:0] RF_WR_ADDR_WB;
  wire   [31:0] ALU_IN1;
  wire   [31:0] RF_OUT2_EXE;
  wire   [31:0] IMM_EXE;
  wire   [31:0] DRAM_IN_EXE;
  wire   [31:0] ALU_IN2;
  wire   [31:0] ALU_OUT;
  wire   [31:0] MULT_OUT;
  wire   [4:0] RF_WR_ADDR_MEM;
  wire   [31:0] LMD_out;
  wire   [31:0] NPC_WB;
  wire   [31:0] ALU_OUT_WB;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37;
  assign \IRAM_ADDR[4]_BAR  = IRAM_ADDR[4];
  assign \IRAM_ADDR[3]_BAR  = IRAM_ADDR[3];
  assign misprediction_BAR = misprediction;

  reg_N32_0 PC ( .D(PC_IN), .EN(\control_from_HDU[PC_EN] ), .CLK(CLK), .RST(
        RST), .\Q[31] (IRAM_ADDR[31]), .\Q[30] (IRAM_ADDR[30]), .\Q[29] (
        IRAM_ADDR[29]), .\Q[28] (IRAM_ADDR[28]), .\Q[27] (IRAM_ADDR[27]), 
        .\Q[26] (IRAM_ADDR[26]), .\Q[25] (IRAM_ADDR[25]), .\Q[24] (
        IRAM_ADDR[24]), .\Q[23] (IRAM_ADDR[23]), .\Q[22] (IRAM_ADDR[22]), 
        .\Q[21] (IRAM_ADDR[21]), .\Q[20] (IRAM_ADDR[20]), .\Q[19] (
        IRAM_ADDR[19]), .\Q[18] (IRAM_ADDR[18]), .\Q[17] (IRAM_ADDR[17]), 
        .\Q[16] (IRAM_ADDR[16]), .\Q[15] (IRAM_ADDR[15]), .\Q[14] (
        IRAM_ADDR[14]), .\Q[13] (IRAM_ADDR[13]), .\Q[12] (IRAM_ADDR[12]), 
        .\Q[11] (IRAM_ADDR[11]), .\Q[10] (IRAM_ADDR[10]), .\Q[9] (IRAM_ADDR[9]), .\Q[8] (IRAM_ADDR[8]), .\Q[7] (IRAM_ADDR[7]), .\Q[6] (IRAM_ADDR[6]), 
        .\Q[5] (IRAM_ADDR[5]), .\Q[1] (IRAM_ADDR[1]), .\Q[0] (IRAM_ADDR[0]), 
        .\Q[3]_BAR (IRAM_ADDR[3]), .\Q[2] (IRAM_ADDR[2]), .\Q[4]_BAR (
        IRAM_ADDR[4]) );
  RCA_N32 ADDER_PC ( .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0}), 
        .Ci(1'b0), .\A[31] (IRAM_ADDR[31]), .\A[30] (IRAM_ADDR[30]), .\A[29] (
        IRAM_ADDR[29]), .\A[28] (IRAM_ADDR[28]), .\A[27] (IRAM_ADDR[27]), 
        .\A[26] (IRAM_ADDR[26]), .\A[25] (IRAM_ADDR[25]), .\A[24] (
        IRAM_ADDR[24]), .\A[23] (IRAM_ADDR[23]), .\A[22] (IRAM_ADDR[22]), 
        .\A[21] (IRAM_ADDR[21]), .\A[20] (IRAM_ADDR[20]), .\A[19] (
        IRAM_ADDR[19]), .\A[18] (IRAM_ADDR[18]), .\A[17] (IRAM_ADDR[17]), 
        .\A[16] (IRAM_ADDR[16]), .\A[15] (IRAM_ADDR[15]), .\A[14] (
        IRAM_ADDR[14]), .\A[13] (IRAM_ADDR[13]), .\A[12] (IRAM_ADDR[12]), 
        .\A[11] (IRAM_ADDR[11]), .\A[10] (IRAM_ADDR[10]), .\A[9] (IRAM_ADDR[9]), .\A[8] (IRAM_ADDR[8]), .\A[7] (IRAM_ADDR[7]), .\A[6] (IRAM_ADDR[6]), 
        .\A[5] (IRAM_ADDR[5]), .\A[1] (IRAM_ADDR[1]), .\A[0] (IRAM_ADDR[0]), 
        .\A[3]_BAR (IRAM_ADDR[3]), .\A[2] (IRAM_ADDR[2]), .\S[31] (NPC[31]), 
        .\S[30] (NPC[30]), .\S[29] (NPC[29]), .\S[28] (NPC[28]), .\S[27] (
        NPC[27]), .\S[26] (NPC[26]), .\S[25] (NPC[25]), .\S[24] (NPC[24]), 
        .\S[23] (NPC[23]), .\S[22] (NPC[22]), .\S[21] (NPC[21]), .\S[20] (
        NPC[20]), .\S[19] (NPC[19]), .\S[18] (NPC[18]), .\S[17] (NPC[17]), 
        .\S[16] (NPC[16]), .\S[15] (NPC[15]), .\S[14] (NPC[14]), .\S[13] (
        NPC[13]), .\S[12] (NPC[12]), .\S[11] (NPC[11]), .\S[10] (NPC[10]), 
        .\S[9] (NPC[9]), .\S[8] (NPC[8]), .\S[7] (NPC[7]), .\S[6] (NPC[6]), 
        .\S[5] (NPC[5]), .\S[4] (NPC[4]), .\S[3] (NPC[3]), .\S[2]_BAR (NPC[2]), 
        .\S[1] (NPC[1]), .\S[0] (NPC[0]), .\A[4]_BAR (IRAM_ADDR[4]) );
  BPU_TAG_FIELD_SIZE8_SET_FIELD_SIZE3_LINES_PER_SET4 BPU_instance ( .clk(CLK), 
        .rst(RST), .instr_fetch({IRAM_OUT[31:27], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .pc_out(
        PC_IN), .actual_addr({actual_addr[31:23], n10, actual_addr[21], n11, 
        actual_addr[19:0]}), .ID_EN(\control_from_HDU[ID_EN] ), .IF_EN(
        \control_from_HDU[IF_EN] ), .\pc_fetch[31] (1'b0), .\pc_fetch[30] (
        1'b0), .\pc_fetch[29] (1'b0), .\pc_fetch[28] (1'b0), .\pc_fetch[27] (
        1'b0), .\pc_fetch[26] (1'b0), .\pc_fetch[25] (1'b0), .\pc_fetch[24] (
        1'b0), .\pc_fetch[23] (1'b0), .\pc_fetch[22] (1'b0), .\pc_fetch[21] (
        1'b0), .\pc_fetch[20] (1'b0), .\pc_fetch[19] (1'b0), .\pc_fetch[18] (
        1'b0), .\pc_fetch[17] (1'b0), .\pc_fetch[16] (1'b0), .\pc_fetch[15] (
        1'b0), .\pc_fetch[14] (1'b0), .\pc_fetch[13] (1'b0), .\pc_fetch[12] (
        IRAM_ADDR[12]), .\pc_fetch[11] (IRAM_ADDR[11]), .\pc_fetch[10] (
        IRAM_ADDR[10]), .\pc_fetch[9] (IRAM_ADDR[9]), .\pc_fetch[8] (
        IRAM_ADDR[8]), .\pc_fetch[7] (IRAM_ADDR[7]), .\pc_fetch[6] (
        IRAM_ADDR[6]), .\pc_fetch[5] (IRAM_ADDR[5]), .\pc_fetch[1] (1'b0), 
        .\pc_fetch[0] (1'b0), .\pc_fetch[3]_BAR (IRAM_ADDR[3]), 
        .misprediction_BAR(misprediction), .\pc_fetch[2] (IRAM_ADDR[2]), 
        .\pc_in[31] (NPC[31]), .\pc_in[30] (NPC[30]), .\pc_in[29] (NPC[29]), 
        .\pc_in[28] (NPC[28]), .\pc_in[27] (NPC[27]), .\pc_in[26] (NPC[26]), 
        .\pc_in[25] (NPC[25]), .\pc_in[24] (NPC[24]), .\pc_in[23] (NPC[23]), 
        .\pc_in[22] (NPC[22]), .\pc_in[21] (NPC[21]), .\pc_in[20] (NPC[20]), 
        .\pc_in[19] (NPC[19]), .\pc_in[18] (NPC[18]), .\pc_in[17] (NPC[17]), 
        .\pc_in[16] (NPC[16]), .\pc_in[15] (NPC[15]), .\pc_in[14] (NPC[14]), 
        .\pc_in[13] (NPC[13]), .\pc_in[12] (NPC[12]), .\pc_in[11] (NPC[11]), 
        .\pc_in[10] (NPC[10]), .\pc_in[9] (NPC[9]), .\pc_in[8] (NPC[8]), 
        .\pc_in[7] (NPC[7]), .\pc_in[6] (NPC[6]), .\pc_in[5] (NPC[5]), 
        .\pc_in[4] (NPC[4]), .\pc_in[3] (NPC[3]), .\pc_in[2]_BAR (1'b0), 
        .\pc_in[1] (NPC[1]), .\pc_in[0] (NPC[0]), .\pc_fetch[4]_BAR (
        IRAM_ADDR[4]) );
  reg_N32_12 REG_NPC_IF ( .Q(NPC_ID), .EN(\control_from_HDU[IF_EN] ), .CLK(CLK), .RST(RST), .\D[31] (NPC[31]), .\D[30] (NPC[30]), .\D[29] (NPC[29]), 
        .\D[28] (NPC[28]), .\D[27] (NPC[27]), .\D[26] (NPC[26]), .\D[25] (
        NPC[25]), .\D[24] (NPC[24]), .\D[23] (NPC[23]), .\D[22] (NPC[22]), 
        .\D[21] (NPC[21]), .\D[20] (NPC[20]), .\D[19] (NPC[19]), .\D[18] (
        NPC[18]), .\D[17] (NPC[17]), .\D[16] (NPC[16]), .\D[15] (NPC[15]), 
        .\D[14] (NPC[14]), .\D[13] (NPC[13]), .\D[12] (NPC[12]), .\D[11] (
        NPC[11]), .\D[10] (NPC[10]), .\D[9] (NPC[9]), .\D[8] (NPC[8]), 
        .\D[7] (NPC[7]), .\D[6] (NPC[6]), .\D[5] (NPC[5]), .\D[4] (NPC[4]), 
        .\D[3] (NPC[3]), .\D[2]_BAR (NPC[2]), .\D[1] (NPC[1]), .\D[0] (NPC[0])
         );
  reg_N32_11 IR ( .D({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, IRAM_OUT[25:0]}), 
        .Q({SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, IR_out}), .EN(
        \control_from_HDU[IF_EN] ), .CLK(CLK), .RST(RST) );
  MUX_2to1_N32_0 MUX_BRANCH ( .IN0({n53, RF_OUT1_fw[30:1], n54}), .IN1(
        ADDER_BRANCH_out), .SEL(\control_from_CU[ID][MUX_BRANCH_SEL] ), .Y(
        NPC_BRANCH) );
  ADDER_P4_N_BIT32_0 ADDER_BRANCH ( .A(NPC_ID), .B({n52, n51, n50, n49, n48, 
        n47, n46, IMM_ID[24:0]}), .add_sub(1'b0), .SUM(ADDER_BRANCH_out) );
  branch_comp_N32 branch_comp_instance ( .BRANCH_COND({
        \control_from_CU[ID][BRANCH_COND][1] , 
        \control_from_CU[ID][BRANCH_COND][0] }), .DATA_IN(RF_OUT1_fw), 
        .BRANCH_IS_TAKEN(branch_is_taken) );
  MUX_2to1_N32_9 MUX_actual_addr ( .IN0(NPC_ID), .IN1(NPC_BRANCH), .SEL(
        branch_is_taken), .Y({actual_addr[31:23], n10, actual_addr[21], n11, 
        actual_addr[19:0]}) );
  MUX_8to1_N32_0 MUX_RF_OUT1_fw ( .IN0(RF_OUT1), .IN1(ALU_OUT_EXE), .IN2(
        DRAM_ADDR), .IN3(LMD_in), .IN4({n16, n21, n37, n39, n25, n33, n42, n34, 
        n14, n27, n31, n29, n32, n36, n41, n35, n40, n12, n28, n43, n38, n22, 
        n24, n17, n19, n20, n18, n23, n30, n15, n26, n13}), .IN5(NPC_MEM), 
        .IN6(NPC_EXE), .IN7({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .SEL({\control_from_FU[MUX_RF_OUT1_SEL][2] , 
        \control_from_FU[MUX_RF_OUT1_SEL][1] , 
        \control_from_FU[MUX_RF_OUT1_SEL][0] }), .Y(RF_OUT1_fw) );
  MUX_8to1_N32_3 MUX_RF_OUT2_fw ( .IN0(RF_OUT2), .IN1({n55, ALU_OUT_EXE[30:8], 
        n8, ALU_OUT_EXE[6:1], n56}), .IN2(DRAM_ADDR), .IN3(LMD_in), .IN4({n16, 
        n21, n37, n39, n25, n33, n42, n34, n14, n27, n31, n29, n32, n36, n41, 
        n35, n40, n12, n28, n43, n38, n22, n24, n17, n19, n20, n18, n23, n30, 
        n15, n26, n13}), .IN5(NPC_MEM), .IN6(NPC_EXE), .IN7({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .SEL({
        \control_from_FU[MUX_RF_OUT2_SEL][2] , 
        \control_from_FU[MUX_RF_OUT2_SEL][1] , 
        \control_from_FU[MUX_RF_OUT2_SEL][0] }), .Y(RF_OUT2_fw) );
  reg_N32_10 REG_NPC_ID ( .D(NPC_ID), .Q(NPC_EXE), .EN(
        \control_from_HDU[ID_EN] ), .CLK(CLK), .RST(RST) );
  MUX_4to1_N5 MUX_RF_WR_ADDR ( .IN0(IR_out[20:16]), .IN1(IR_out[15:11]), .IN2(
        {1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .IN3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL({\control_from_CU[ID][MUX_RF_WR_ADDR_SEL][1] , 
        \control_from_CU[ID][MUX_RF_WR_ADDR_SEL][0] }), .Y(RF_WR_ADDR_ID) );
  reg_N5_0 REG_RF_WR_ADDR_ID ( .D(RF_WR_ADDR_ID), .Q(RF_WR_ADDR_EXE), .EN(
        \control_from_HDU[ID_EN] ), .CLK(CLK), .RST(RST) );
  RF_N_bit32_N_reg32 RF_instance ( .CLK(CLK), .RST(RST), .WR_EN(
        \control_from_CU[WB][RF_WR_EN] ), .ADD_WR(RF_WR_ADDR_WB), .ADD_RD1(
        IR_out[25:21]), .ADD_RD2(IR_out[20:16]), .DATA_IN({n16, n21, n37, n39, 
        n25, n33, n42, n34, n14, n27, n31, n29, n32, n36, n41, n35, n40, n12, 
        n28, n43, n38, n22, n24, n17, n19, n20, n18, n23, n30, n15, n26, n13}), 
        .OUT1(RF_OUT1), .OUT2(RF_OUT2) );
  reg_N32_9 REG_RF_OUT1 ( .D({n53, RF_OUT1_fw[30:1], n54}), .EN(
        \control_from_HDU[ID_EN] ), .CLK(CLK), .RST(RST), .\Q[31] (ALU_IN1[31]), .\Q[30] (ALU_IN1[30]), .\Q[29] (ALU_IN1[29]), .\Q[28] (ALU_IN1[28]), 
        .\Q[27] (ALU_IN1[27]), .\Q[26] (ALU_IN1[26]), .\Q[25] (ALU_IN1[25]), 
        .\Q[24] (ALU_IN1[24]), .\Q[23] (ALU_IN1[23]), .\Q[22] (ALU_IN1[22]), 
        .\Q[21] (ALU_IN1[21]), .\Q[20]_BAR (ALU_IN1[20]), .\Q[17] (ALU_IN1[17]), .\Q[15] (ALU_IN1[15]), .\Q[11] (ALU_IN1[11]), .\Q[10] (ALU_IN1[10]), 
        .\Q[9] (ALU_IN1[9]), .\Q[8] (ALU_IN1[8]), .\Q[7] (ALU_IN1[7]), 
        .\Q[6] (ALU_IN1[6]), .\Q[5] (ALU_IN1[5]), .\Q[4] (ALU_IN1[4]), 
        .\Q[3] (ALU_IN1[3]), .\Q[2] (ALU_IN1[2]), .\Q[1] (ALU_IN1[1]), 
        .\Q[0] (ALU_IN1[0]), .\Q[19]_BAR (ALU_IN1[19]), .\Q[18]_BAR (
        ALU_IN1[18]), .\Q[16]_BAR (ALU_IN1[16]), .\Q[14]_BAR (ALU_IN1[14]), 
        .\Q[13]_BAR (ALU_IN1[13]), .\Q[12]_BAR (ALU_IN1[12]) );
  reg_N32_8 REG_RF_OUT2 ( .D(RF_OUT2_fw), .Q(RF_OUT2_EXE), .EN(
        \control_from_HDU[ID_EN] ), .CLK(CLK), .RST(RST) );
  MUX_2to1_N32_8 MUX_IMM_EXT ( .IN0({IR_out[15], IR_out[15], IR_out[15], 
        IR_out[15], IR_out[15], IR_out[15], IR_out[15], IR_out[15], IR_out[15], 
        IR_out[15], IR_out[15], IR_out[15], IR_out[15], IR_out[15], IR_out[15], 
        IR_out[15], IR_out[15:0]}), .IN1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        IR_out[25:16], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .SEL(
        \control_from_CU[ID][MUX_IMM_EXT_SEL] ), .Y({n52, n51, n50, n49, n48, 
        n47, n46, IMM_ID[24:0]}) );
  reg_N32_7 REG_IMM ( .D({n52, n51, n50, n49, n48, n47, n46, IMM_ID[24:0]}), 
        .Q(IMM_EXE), .EN(\control_from_HDU[ID_EN] ), .CLK(CLK), .RST(RST) );
  MUX_2to1_N32_7 MUX_DRAM_IN_fw ( .IN0(RF_OUT2_EXE), .IN1(LMD_in), .SEL(
        \control_from_FU[MUX_DRAM_IN_SEL] ), .Y(DRAM_IN_EXE) );
  MUX_2to1_N32_6 MUX_ALU_IN2 ( .IN0(RF_OUT2_EXE), .IN1(IMM_EXE), .SEL(
        \control_from_CU[EXE][MUX_ALU_IN2_SEL] ), .Y({ALU_IN2[31:26], n44, 
        ALU_IN2[24:10], n45, ALU_IN2[8:0]}) );
  ALU_N32 ALU_instance ( .FUNC({\control_from_CU[EXE][ALU_OP][4] , 
        \control_from_CU[EXE][ALU_OP][3] , \control_from_CU[EXE][ALU_OP][2] , 
        \control_from_CU[EXE][ALU_OP][1] , \control_from_CU[EXE][ALU_OP][0] }), 
        .DATA1({ALU_IN1[31:21], n7, n6, n5, ALU_IN1[17], n4, ALU_IN1[15], n3, 
        n2, n1, ALU_IN1[11:4], n57, n155, n157, n156}), .DATA2({ALU_IN2[31:26], 
        n44, ALU_IN2[24:11], n58, n45, ALU_IN2[8:3], n9, n59, ALU_IN2[0]}), 
        .OUT_ALU(ALU_OUT) );
  boothmul_4stage_N32 MULT ( .A({ALU_IN1[31:21], n7, n6, n5, ALU_IN1[17], n4, 
        ALU_IN1[15], n3, n2, n1, ALU_IN1[11:0]}), .B({ALU_IN2[31:26], n44, 
        ALU_IN2[24:10], n45, ALU_IN2[8:0]}), .EN(
        \control_from_CU[EXE][MULT_EN] ), .CLK(CLK), .RST(RST), .P({
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, MULT_OUT}) );
  MUX_2to1_N32_5 MUX_MULT ( .IN0(ALU_OUT), .IN1(MULT_OUT), .SEL(
        \control_from_CU[EXE][MUX_MULT_SEL] ), .Y(ALU_OUT_EXE) );
  reg_N32_6 REG_ALU_OUT_EXE ( .D({n55, ALU_OUT_EXE[30:8], n8, ALU_OUT_EXE[6:1], 
        n56}), .Q(DRAM_ADDR), .EN(\control_from_HDU[EXE_EN] ), .CLK(CLK), 
        .RST(RST) );
  reg_N32_5 REG_NPC_EXE ( .D(NPC_EXE), .Q(NPC_MEM), .EN(
        \control_from_HDU[EXE_EN] ), .CLK(CLK), .RST(RST) );
  reg_N32_4 REG_DRAM_IN ( .D(DRAM_IN_EXE), .Q(DRAM_IN), .EN(
        \control_from_HDU[EXE_EN] ), .CLK(CLK), .RST(RST) );
  reg_N5_2 REG_RF_WR_ADDR_EXE ( .D(RF_WR_ADDR_EXE), .Q(RF_WR_ADDR_MEM), .EN(
        \control_from_HDU[EXE_EN] ), .CLK(CLK), .RST(RST) );
  MUX_8to1_N32_2 MUX_DRAM_OUT_EXT ( .IN0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, DRAM_OUT[7], 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .IN1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .IN2({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, DRAM_OUT[15], 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .IN3({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN4({DRAM_OUT[31:16], 1'b0, DRAM_OUT[14:8], 1'b0, DRAM_OUT[6:0]}), .IN5({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN6({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .IN7({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .SEL({
        \control_from_CU[MEM][MUX_DRAM_OUT_EXT_SEL][2] , 
        \control_from_CU[MEM][MUX_DRAM_OUT_EXT_SEL][1] , 
        \control_from_CU[MEM][MUX_DRAM_OUT_EXT_SEL][0] }), .Y(LMD_in) );
  reg_N32_3 LMD ( .D(LMD_in), .Q(LMD_out), .EN(1'b1), .CLK(CLK), .RST(RST) );
  reg_N32_2 REG_NPC_MEM ( .D(NPC_MEM), .Q(NPC_WB), .EN(1'b1), .CLK(CLK), .RST(
        RST) );
  reg_N32_1 REG_ALU_OUT_MEM ( .D(DRAM_ADDR), .Q(ALU_OUT_WB), .EN(1'b1), .CLK(
        CLK), .RST(RST) );
  reg_N5_1 REG_RF_WR_ADDR_MEM ( .D(RF_WR_ADDR_MEM), .Q(RF_WR_ADDR_WB), .EN(
        1'b1), .CLK(CLK), .RST(RST) );
  MUX_4to1_N32 MUX_WB ( .IN0(NPC_WB), .IN1(LMD_out), .IN2(ALU_OUT_WB), .IN3({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .SEL({
        \control_from_CU[WB][MUX_WB_SEL][1] , 
        \control_from_CU[WB][MUX_WB_SEL][0] }), .Y({n16, n21, n37, n39, n25, 
        n33, n42, n34, n14, n27, n31, n29, n32, n36, n41, n35, n40, n12, n28, 
        n43, n38, n22, n24, n17, n19, n20, n18, n23, n30, n15, n26, n13}) );
  INV_X2 U4 ( .A(ALU_IN1[12]), .ZN(n1) );
  INV_X2 U5 ( .A(ALU_IN1[13]), .ZN(n2) );
  INV_X2 U6 ( .A(ALU_IN1[14]), .ZN(n3) );
  INV_X2 U7 ( .A(ALU_IN1[16]), .ZN(n4) );
  INV_X2 U8 ( .A(ALU_IN1[18]), .ZN(n5) );
  INV_X2 U9 ( .A(ALU_IN1[19]), .ZN(n6) );
  INV_X2 U10 ( .A(ALU_IN1[20]), .ZN(n7) );
  BUF_X1 U11 ( .A(ALU_OUT_EXE[7]), .Z(n8) );
  BUF_X1 U12 ( .A(ALU_IN2[2]), .Z(n9) );
  BUF_X1 U13 ( .A(RF_OUT1_fw[31]), .Z(n53) );
  BUF_X1 U14 ( .A(ALU_OUT_EXE[31]), .Z(n55) );
  BUF_X1 U15 ( .A(ALU_IN2[1]), .Z(n59) );
  BUF_X1 U16 ( .A(ALU_IN2[10]), .Z(n58) );
  BUF_X1 U17 ( .A(ALU_IN1[3]), .Z(n57) );
  BUF_X1 U18 ( .A(ALU_IN1[2]), .Z(n155) );
  BUF_X1 U19 ( .A(ALU_IN1[1]), .Z(n157) );
  BUF_X1 U20 ( .A(RF_OUT1_fw[0]), .Z(n54) );
  BUF_X1 U21 ( .A(ALU_OUT_EXE[0]), .Z(n56) );
  BUF_X1 U22 ( .A(ALU_IN1[0]), .Z(n156) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_DLX_BPU_TAG_FIELD_SIZE8_BPU_SET_FIELD_SIZE3_BPU_LINES_PER_SET4_5 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18716, net18718, net18720, net18721, net18724, net18727;
  assign net18716 = EN;
  assign net18718 = CLK;
  assign ENCLK = net18720;
  assign net18727 = TE;

  DLL_X1 latch ( .D(net18721), .GN(net18718), .Q(net18724) );
  AND2_X1 main_gate ( .A1(net18724), .A2(net18718), .ZN(net18720) );
  OR2_X1 test_or ( .A1(net18716), .A2(net18727), .ZN(net18721) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_DLX_BPU_TAG_FIELD_SIZE8_BPU_SET_FIELD_SIZE3_BPU_LINES_PER_SET4_4 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18716, net18718, net18720, net18721, net18724, net18727;
  assign net18716 = EN;
  assign net18718 = CLK;
  assign ENCLK = net18720;
  assign net18727 = TE;

  DLL_X1 latch ( .D(net18721), .GN(net18718), .Q(net18724) );
  AND2_X1 main_gate ( .A1(net18724), .A2(net18718), .ZN(net18720) );
  OR2_X1 test_or ( .A1(net18716), .A2(net18727), .ZN(net18721) );
endmodule



    module SNPS_CLOCK_GATE_HIGH_DLX_BPU_TAG_FIELD_SIZE8_BPU_SET_FIELD_SIZE3_BPU_LINES_PER_SET4_3 ( 
        CLK, EN, ENCLK, TE );
  input CLK, EN, TE;
  output ENCLK;
  wire   net18716, net18718, net18720, net18721, net18724, net18727;
  assign net18716 = EN;
  assign net18718 = CLK;
  assign ENCLK = net18720;
  assign net18727 = TE;

  DLL_X1 latch ( .D(net18721), .GN(net18718), .Q(net18724) );
  AND2_X1 main_gate ( .A1(net18724), .A2(net18718), .ZN(net18720) );
  OR2_X1 test_or ( .A1(net18716), .A2(net18727), .ZN(net18721) );
endmodule


module DLX_BPU_TAG_FIELD_SIZE8_BPU_SET_FIELD_SIZE3_BPU_LINES_PER_SET4 ( 
        IRAM_ADDR, IRAM_OUT, DRAM_ADDR, DRAM_IN, DRAM_OUT, .DRAM_WR_EN({
        \DRAM_WR_EN[1] , \DRAM_WR_EN[0] }), CLK, RST );
  output [31:0] IRAM_ADDR;
  input [31:0] IRAM_OUT;
  output [31:0] DRAM_ADDR;
  output [31:0] DRAM_IN;
  input [31:0] DRAM_OUT;
  input CLK, RST;
  output \DRAM_WR_EN[1] , \DRAM_WR_EN[0] ;
  wire   n215, n216, \HDU_OUTS[PC_EN] , \HDU_OUTS[IF_EN] , \HDU_OUTS[ID_EN] ,
         \HDU_OUTS[EXE_EN] , \HDU_OUTS[ID_BUBBLE] , \HDU_OUTS[EXE_BUBBLE] ,
         \HDU_OUTS[MEM_BUBBLE] , N5, N32, N34, N36, N39, N66, N68, N70, N100,
         N102, N104, N134, N136, N138, misprediction,
         \FU_OUTS[MUX_RF_OUT1_SEL][2] , \FU_OUTS[MUX_RF_OUT1_SEL][1] ,
         \FU_OUTS[MUX_RF_OUT1_SEL][0] , \FU_OUTS[MUX_RF_OUT2_SEL][2] ,
         \FU_OUTS[MUX_RF_OUT2_SEL][1] , \FU_OUTS[MUX_RF_OUT2_SEL][0] ,
         \FU_OUTS[MUX_DRAM_IN_SEL] , \CU_OUTS[ID][MUX_BRANCH_SEL] ,
         \CU_OUTS[ID][MUX_IMM_EXT_SEL] , \CU_OUTS[ID][MUX_RF_WR_ADDR_SEL][1] ,
         \CU_OUTS[ID][MUX_RF_WR_ADDR_SEL][0] , \CU_OUTS[ID][BRANCH_COND][1] ,
         \CU_OUTS[ID][BRANCH_COND][0] , \CU_OUTS[EXE][MULT_EN] ,
         \CU_OUTS[EXE][MUX_MULT_SEL] , \CU_OUTS[EXE][ALU_OP][4] ,
         \CU_OUTS[EXE][ALU_OP][3] , \CU_OUTS[EXE][ALU_OP][2] ,
         \CU_OUTS[EXE][ALU_OP][1] , \CU_OUTS[EXE][ALU_OP][0] ,
         \CU_OUTS[MEM][DRAM_WR_EN][1] , \CU_OUTS[MEM][DRAM_WR_EN][0] ,
         \CU_OUTS[MEM][MUX_DRAM_OUT_EXT_SEL][2] ,
         \CU_OUTS[MEM][MUX_DRAM_OUT_EXT_SEL][1] ,
         \CU_OUTS[MEM][MUX_DRAM_OUT_EXT_SEL][0] , \CU_OUTS[WB][MUX_WB_SEL][1] ,
         \CU_OUTS[WB][MUX_WB_SEL][0] , \CU_OUTS[WB][RF_WR_EN] ,
         \CU_OUTS_EXE_atEXE[MULT_EN] , \CU_OUTS_EXE_atEXE[MUX_MULT_SEL] ,
         \CU_OUTS_EXE_atEXE[MUX_ALU_IN2_SEL] , \CU_OUTS_EXE_atEXE[ALU_OP][4] ,
         \CU_OUTS_EXE_atEXE[ALU_OP][3] , \CU_OUTS_EXE_atEXE[ALU_OP][2] ,
         \CU_OUTS_EXE_atEXE[ALU_OP][1] , \CU_OUTS_EXE_atEXE[ALU_OP][0] ,
         \CU_OUTS_MEM_atEXE[DRAM_WR_EN][1] ,
         \CU_OUTS_MEM_atEXE[DRAM_WR_EN][0] , \CU_OUTS_WB_atEXE[RF_WR_EN] ,
         \CU_OUTS_MEM_atMEM[MUX_DRAM_OUT_EXT_SEL][2] ,
         \CU_OUTS_MEM_atMEM[MUX_DRAM_OUT_EXT_SEL][1] ,
         \CU_OUTS_MEM_atMEM[MUX_DRAM_OUT_EXT_SEL][0] ,
         \CU_OUTS_WB_atMEM[RF_WR_EN] , \CU_OUTS_WB_atWB[MUX_WB_SEL][1] ,
         \CU_OUTS_WB_atWB[MUX_WB_SEL][0] , \CU_OUTS_WB_atWB[RF_WR_EN] ,
         net18743, net18748, net18753, n14, n15, n16, n17, n18, n19, n20, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210;
  wire   [1:0] DRAM_WR_EN;
  wire   [31:0] INSTR_ID;
  wire   [31:0] INSTR_EXE;
  wire   [31:0] INSTR_MEM;
  wire   [31:0] INSTR_WB;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  HDU HDU_instance ( .INSTR_ID({INSTR_ID[31:16], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .INSTR_EXE({INSTR_EXE[31:26], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        INSTR_EXE[20:16], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, INSTR_EXE[5:0]}), .HDU_OUTS({\HDU_OUTS[PC_EN] , 
        \HDU_OUTS[IF_EN] , \HDU_OUTS[ID_EN] , \HDU_OUTS[EXE_EN] , 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        \HDU_OUTS[ID_BUBBLE] , \HDU_OUTS[EXE_BUBBLE] , \HDU_OUTS[MEM_BUBBLE] , 
        SYNOPSYS_UNCONNECTED__2}), .clk(CLK), .rst(RST), .misprediction_BAR(
        misprediction) );
  FU FU_instance ( .INSTR_ID({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        INSTR_ID[25:16], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .INSTR_EXE({
        INSTR_EXE[31:26], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, INSTR_EXE[20:11], 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .INSTR_MEM({INSTR_MEM[31], N138, INSTR_MEM[29], N136, INSTR_MEM[27], 
        N134, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, INSTR_MEM[20:11], 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .INSTR_WB({
        INSTR_WB[31:26], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, INSTR_WB[20:11], 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .FU_OUTS({\FU_OUTS[MUX_RF_OUT1_SEL][2] , \FU_OUTS[MUX_RF_OUT1_SEL][1] , 
        \FU_OUTS[MUX_RF_OUT1_SEL][0] , \FU_OUTS[MUX_RF_OUT2_SEL][2] , 
        \FU_OUTS[MUX_RF_OUT2_SEL][1] , \FU_OUTS[MUX_RF_OUT2_SEL][0] , 
        \FU_OUTS[MUX_DRAM_IN_SEL] }) );
  CU CU_instance ( .INSTR_ID({INSTR_ID[31:26], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, INSTR_ID[5:0]}), .CU_OUTS({
        \CU_OUTS[ID][MUX_BRANCH_SEL] , \CU_OUTS[ID][MUX_IMM_EXT_SEL] , 
        \CU_OUTS[ID][MUX_RF_WR_ADDR_SEL][1] , 
        \CU_OUTS[ID][MUX_RF_WR_ADDR_SEL][0] , \CU_OUTS[ID][BRANCH_COND][1] , 
        \CU_OUTS[ID][BRANCH_COND][0] , \CU_OUTS[EXE][MULT_EN] , 
        \CU_OUTS[EXE][MUX_MULT_SEL] , SYNOPSYS_UNCONNECTED__3, 
        \CU_OUTS[EXE][ALU_OP][4] , \CU_OUTS[EXE][ALU_OP][3] , 
        \CU_OUTS[EXE][ALU_OP][2] , \CU_OUTS[EXE][ALU_OP][1] , 
        \CU_OUTS[EXE][ALU_OP][0] , \CU_OUTS[MEM][DRAM_WR_EN][1] , 
        \CU_OUTS[MEM][DRAM_WR_EN][0] , \CU_OUTS[MEM][MUX_DRAM_OUT_EXT_SEL][2] , 
        \CU_OUTS[MEM][MUX_DRAM_OUT_EXT_SEL][1] , 
        \CU_OUTS[MEM][MUX_DRAM_OUT_EXT_SEL][0] , \CU_OUTS[WB][MUX_WB_SEL][1] , 
        \CU_OUTS[WB][MUX_WB_SEL][0] , \CU_OUTS[WB][RF_WR_EN] }) );
  datapath_BPU_TAG_FIELD_SIZE8_BPU_SET_FIELD_SIZE3_BPU_LINES_PER_SET4 datapath_instance ( 
        .IRAM_OUT({IRAM_OUT[31:27], 1'b0, IRAM_OUT[25:0]}), .DRAM_ADDR(
        DRAM_ADDR), .DRAM_IN(DRAM_IN), .DRAM_OUT(DRAM_OUT), .control_from_CU({
        \CU_OUTS[ID][MUX_BRANCH_SEL] , \CU_OUTS[ID][MUX_IMM_EXT_SEL] , 
        \CU_OUTS[ID][MUX_RF_WR_ADDR_SEL][1] , 
        \CU_OUTS[ID][MUX_RF_WR_ADDR_SEL][0] , \CU_OUTS[ID][BRANCH_COND][1] , 
        \CU_OUTS[ID][BRANCH_COND][0] , \CU_OUTS_EXE_atEXE[MULT_EN] , 
        \CU_OUTS_EXE_atEXE[MUX_MULT_SEL] , 
        \CU_OUTS_EXE_atEXE[MUX_ALU_IN2_SEL] , \CU_OUTS_EXE_atEXE[ALU_OP][4] , 
        \CU_OUTS_EXE_atEXE[ALU_OP][3] , \CU_OUTS_EXE_atEXE[ALU_OP][2] , 
        \CU_OUTS_EXE_atEXE[ALU_OP][1] , \CU_OUTS_EXE_atEXE[ALU_OP][0] , 1'b0, 
        1'b0, \CU_OUTS_MEM_atMEM[MUX_DRAM_OUT_EXT_SEL][2] , 
        \CU_OUTS_MEM_atMEM[MUX_DRAM_OUT_EXT_SEL][1] , 
        \CU_OUTS_MEM_atMEM[MUX_DRAM_OUT_EXT_SEL][0] , 
        \CU_OUTS_WB_atWB[MUX_WB_SEL][1] , \CU_OUTS_WB_atWB[MUX_WB_SEL][0] , 
        \CU_OUTS_WB_atWB[RF_WR_EN] }), .control_from_FU({
        \FU_OUTS[MUX_RF_OUT1_SEL][2] , \FU_OUTS[MUX_RF_OUT1_SEL][1] , 
        \FU_OUTS[MUX_RF_OUT1_SEL][0] , \FU_OUTS[MUX_RF_OUT2_SEL][2] , 
        \FU_OUTS[MUX_RF_OUT2_SEL][1] , \FU_OUTS[MUX_RF_OUT2_SEL][0] , 
        \FU_OUTS[MUX_DRAM_IN_SEL] }), .control_from_HDU({\HDU_OUTS[PC_EN] , 
        \HDU_OUTS[IF_EN] , \HDU_OUTS[ID_EN] , \HDU_OUTS[EXE_EN] , 1'b1, 1'b1, 
        1'b0, 1'b0, 1'b0, 1'b0}), .CLK(CLK), .RST(RST), .\IRAM_ADDR[31] (
        IRAM_ADDR[31]), .\IRAM_ADDR[30] (IRAM_ADDR[30]), .\IRAM_ADDR[29] (
        IRAM_ADDR[29]), .\IRAM_ADDR[28] (IRAM_ADDR[28]), .\IRAM_ADDR[27] (
        IRAM_ADDR[27]), .\IRAM_ADDR[26] (IRAM_ADDR[26]), .\IRAM_ADDR[25] (
        IRAM_ADDR[25]), .\IRAM_ADDR[24] (IRAM_ADDR[24]), .\IRAM_ADDR[23] (
        IRAM_ADDR[23]), .\IRAM_ADDR[22] (IRAM_ADDR[22]), .\IRAM_ADDR[21] (
        IRAM_ADDR[21]), .\IRAM_ADDR[20] (IRAM_ADDR[20]), .\IRAM_ADDR[19] (
        IRAM_ADDR[19]), .\IRAM_ADDR[18] (IRAM_ADDR[18]), .\IRAM_ADDR[17] (
        IRAM_ADDR[17]), .\IRAM_ADDR[16] (IRAM_ADDR[16]), .\IRAM_ADDR[15] (
        IRAM_ADDR[15]), .\IRAM_ADDR[14] (IRAM_ADDR[14]), .\IRAM_ADDR[13] (
        IRAM_ADDR[13]), .\IRAM_ADDR[12] (IRAM_ADDR[12]), .\IRAM_ADDR[11] (
        IRAM_ADDR[11]), .\IRAM_ADDR[10] (IRAM_ADDR[10]), .\IRAM_ADDR[9] (
        IRAM_ADDR[9]), .\IRAM_ADDR[8] (IRAM_ADDR[8]), .\IRAM_ADDR[7] (
        IRAM_ADDR[7]), .\IRAM_ADDR[6] (IRAM_ADDR[6]), .\IRAM_ADDR[5] (
        IRAM_ADDR[5]), .\IRAM_ADDR[1] (IRAM_ADDR[1]), .\IRAM_ADDR[0] (
        IRAM_ADDR[0]), .\IRAM_ADDR[3]_BAR (n216), .misprediction_BAR(
        misprediction), .\IRAM_ADDR[2] (IRAM_ADDR[2]), .\IRAM_ADDR[4]_BAR (
        n215) );
  SNPS_CLOCK_GATE_HIGH_DLX_BPU_TAG_FIELD_SIZE8_BPU_SET_FIELD_SIZE3_BPU_LINES_PER_SET4_5 clk_gate_INSTR_ID_reg ( 
        .CLK(CLK), .EN(N5), .ENCLK(net18743), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_DLX_BPU_TAG_FIELD_SIZE8_BPU_SET_FIELD_SIZE3_BPU_LINES_PER_SET4_4 clk_gate_INSTR_EXE_reg ( 
        .CLK(CLK), .EN(N39), .ENCLK(net18748), .TE(1'b0) );
  SNPS_CLOCK_GATE_HIGH_DLX_BPU_TAG_FIELD_SIZE8_BPU_SET_FIELD_SIZE3_BPU_LINES_PER_SET4_3 clk_gate_INSTR_EXE_reg_0 ( 
        .CLK(CLK), .EN(N39), .ENCLK(net18753), .TE(1'b0) );
  DFFS_X1 \INSTR_ID_reg[30]  ( .D(N36), .CK(net18743), .SN(RST), .Q(
        INSTR_ID[30]) );
  DFFS_X1 \INSTR_EXE_reg[30]  ( .D(N70), .CK(net18748), .SN(RST), .Q(
        INSTR_EXE[30]) );
  DFFS_X1 \INSTR_MEM_reg[30]  ( .D(N104), .CK(CLK), .SN(RST), .Q(N138) );
  DFFS_X1 \INSTR_WB_reg[30]  ( .D(N138), .CK(CLK), .SN(RST), .Q(INSTR_WB[30])
         );
  DFFS_X1 \INSTR_ID_reg[28]  ( .D(N34), .CK(net18743), .SN(RST), .Q(
        INSTR_ID[28]) );
  DFFS_X1 \INSTR_EXE_reg[28]  ( .D(N68), .CK(net18748), .SN(RST), .Q(
        INSTR_EXE[28]) );
  DFFS_X1 \INSTR_MEM_reg[28]  ( .D(N102), .CK(CLK), .SN(RST), .Q(N136) );
  DFFS_X1 \INSTR_WB_reg[28]  ( .D(N136), .CK(CLK), .SN(RST), .Q(INSTR_WB[28])
         );
  DFFS_X1 \INSTR_ID_reg[26]  ( .D(N32), .CK(net18743), .SN(RST), .Q(
        INSTR_ID[26]) );
  DFFS_X1 \INSTR_EXE_reg[26]  ( .D(N66), .CK(net18748), .SN(RST), .Q(
        INSTR_EXE[26]) );
  DFFS_X1 \INSTR_MEM_reg[26]  ( .D(N100), .CK(CLK), .SN(RST), .Q(N134) );
  DFFS_X1 \INSTR_WB_reg[26]  ( .D(N134), .CK(CLK), .SN(RST), .Q(INSTR_WB[26])
         );
  DFF_X1 \CU_OUTS_WB_atEXE_reg[MUX_WB_SEL][0]  ( .D(
        \CU_OUTS[WB][MUX_WB_SEL][0] ), .CK(net18753), .QN(n20) );
  DFF_X1 \CU_OUTS_WB_atMEM_reg[MUX_WB_SEL][0]  ( .D(n20), .CK(CLK), .Q(n19) );
  DFF_X1 \CU_OUTS_WB_atWB_reg[MUX_WB_SEL][0]  ( .D(n19), .CK(CLK), .QN(
        \CU_OUTS_WB_atWB[MUX_WB_SEL][0] ) );
  DFF_X1 \CU_OUTS_WB_atEXE_reg[MUX_WB_SEL][1]  ( .D(
        \CU_OUTS[WB][MUX_WB_SEL][1] ), .CK(net18753), .QN(n18) );
  DFF_X1 \CU_OUTS_WB_atMEM_reg[MUX_WB_SEL][1]  ( .D(n18), .CK(CLK), .Q(n17) );
  DFF_X1 \CU_OUTS_WB_atWB_reg[MUX_WB_SEL][1]  ( .D(n17), .CK(CLK), .QN(
        \CU_OUTS_WB_atWB[MUX_WB_SEL][1] ) );
  DFF_X1 \CU_OUTS_MEM_atEXE_reg[MUX_DRAM_OUT_EXT_SEL][0]  ( .D(
        \CU_OUTS[MEM][MUX_DRAM_OUT_EXT_SEL][0] ), .CK(net18753), .QN(n16) );
  DFF_X1 \CU_OUTS_MEM_atMEM_reg[MUX_DRAM_OUT_EXT_SEL][0]  ( .D(n16), .CK(CLK), 
        .QN(\CU_OUTS_MEM_atMEM[MUX_DRAM_OUT_EXT_SEL][0] ) );
  DFF_X1 \CU_OUTS_MEM_atEXE_reg[MUX_DRAM_OUT_EXT_SEL][1]  ( .D(
        \CU_OUTS[MEM][MUX_DRAM_OUT_EXT_SEL][1] ), .CK(net18753), .QN(n15) );
  DFF_X1 \CU_OUTS_MEM_atMEM_reg[MUX_DRAM_OUT_EXT_SEL][1]  ( .D(n15), .CK(CLK), 
        .QN(\CU_OUTS_MEM_atMEM[MUX_DRAM_OUT_EXT_SEL][1] ) );
  DFF_X1 \CU_OUTS_MEM_atEXE_reg[MUX_DRAM_OUT_EXT_SEL][2]  ( .D(
        \CU_OUTS[MEM][MUX_DRAM_OUT_EXT_SEL][2] ), .CK(net18753), .QN(n14) );
  DFF_X1 \CU_OUTS_MEM_atMEM_reg[MUX_DRAM_OUT_EXT_SEL][2]  ( .D(n14), .CK(CLK), 
        .QN(\CU_OUTS_MEM_atMEM[MUX_DRAM_OUT_EXT_SEL][2] ) );
  DFF_X1 \CU_OUTS_EXE_atEXE_reg[MUX_MULT_SEL]  ( .D(
        \CU_OUTS[EXE][MUX_MULT_SEL] ), .CK(net18753), .Q(
        \CU_OUTS_EXE_atEXE[MUX_MULT_SEL] ) );
  DFFS_X1 \CU_OUTS_EXE_atEXE_reg[ALU_OP][3]  ( .D(n209), .CK(net18753), .SN(
        RST), .QN(\CU_OUTS_EXE_atEXE[ALU_OP][3] ) );
  DFFS_X1 \CU_OUTS_EXE_atEXE_reg[ALU_OP][2]  ( .D(n206), .CK(net18753), .SN(
        RST), .QN(\CU_OUTS_EXE_atEXE[ALU_OP][2] ) );
  DFFS_X1 \CU_OUTS_EXE_atEXE_reg[ALU_OP][1]  ( .D(n208), .CK(net18753), .SN(
        RST), .QN(\CU_OUTS_EXE_atEXE[ALU_OP][1] ) );
  DFFS_X1 \CU_OUTS_EXE_atEXE_reg[ALU_OP][0]  ( .D(n207), .CK(net18753), .SN(
        RST), .QN(\CU_OUTS_EXE_atEXE[ALU_OP][0] ) );
  DFF_X1 \CU_OUTS_EXE_atEXE_reg[MUX_ALU_IN2_SEL]  ( .D(
        \CU_OUTS[ID][MUX_RF_WR_ADDR_SEL][0] ), .CK(net18753), .QN(
        \CU_OUTS_EXE_atEXE[MUX_ALU_IN2_SEL] ) );
  DFFR_X1 \CU_OUTS_WB_atWB_reg[RF_WR_EN]  ( .D(\CU_OUTS_WB_atMEM[RF_WR_EN] ), 
        .CK(CLK), .RN(RST), .Q(\CU_OUTS_WB_atWB[RF_WR_EN] ) );
  DFFR_X1 \INSTR_WB_reg[20]  ( .D(INSTR_MEM[20]), .CK(CLK), .RN(RST), .Q(
        INSTR_WB[20]) );
  DFFR_X1 \INSTR_WB_reg[19]  ( .D(INSTR_MEM[19]), .CK(CLK), .RN(RST), .Q(
        INSTR_WB[19]) );
  DFFR_X1 \INSTR_WB_reg[18]  ( .D(INSTR_MEM[18]), .CK(CLK), .RN(RST), .Q(
        INSTR_WB[18]) );
  DFFR_X1 \INSTR_WB_reg[17]  ( .D(INSTR_MEM[17]), .CK(CLK), .RN(RST), .Q(
        INSTR_WB[17]) );
  DFFR_X1 \INSTR_WB_reg[16]  ( .D(INSTR_MEM[16]), .CK(CLK), .RN(RST), .Q(
        INSTR_WB[16]) );
  DFFR_X1 \INSTR_WB_reg[15]  ( .D(INSTR_MEM[15]), .CK(CLK), .RN(RST), .Q(
        INSTR_WB[15]) );
  DFFR_X1 \INSTR_WB_reg[14]  ( .D(INSTR_MEM[14]), .CK(CLK), .RN(RST), .Q(
        INSTR_WB[14]) );
  DFFR_X1 \INSTR_WB_reg[13]  ( .D(INSTR_MEM[13]), .CK(CLK), .RN(RST), .Q(
        INSTR_WB[13]) );
  DFFR_X1 \INSTR_WB_reg[12]  ( .D(INSTR_MEM[12]), .CK(CLK), .RN(RST), .Q(
        INSTR_WB[12]) );
  DFFR_X1 \INSTR_WB_reg[11]  ( .D(INSTR_MEM[11]), .CK(CLK), .RN(RST), .Q(
        INSTR_WB[11]) );
  DFFR_X1 \INSTR_WB_reg[29]  ( .D(INSTR_MEM[29]), .CK(CLK), .RN(RST), .Q(
        INSTR_WB[29]) );
  DFFR_X1 \INSTR_WB_reg[27]  ( .D(INSTR_MEM[27]), .CK(CLK), .RN(RST), .Q(
        INSTR_WB[27]) );
  DFFR_X1 \INSTR_WB_reg[31]  ( .D(INSTR_MEM[31]), .CK(CLK), .RN(RST), .Q(
        INSTR_WB[31]) );
  DFFR_X1 \INSTR_MEM_reg[31]  ( .D(n203), .CK(CLK), .RN(RST), .Q(INSTR_MEM[31]) );
  DFFR_X1 \INSTR_MEM_reg[29]  ( .D(n202), .CK(CLK), .RN(RST), .Q(INSTR_MEM[29]) );
  DFFR_X1 \INSTR_MEM_reg[27]  ( .D(n201), .CK(CLK), .RN(RST), .Q(INSTR_MEM[27]) );
  DFFR_X1 \INSTR_MEM_reg[20]  ( .D(n200), .CK(CLK), .RN(RST), .Q(INSTR_MEM[20]) );
  DFFR_X1 \INSTR_MEM_reg[19]  ( .D(n199), .CK(CLK), .RN(RST), .Q(INSTR_MEM[19]) );
  DFFR_X1 \INSTR_MEM_reg[18]  ( .D(n198), .CK(CLK), .RN(RST), .Q(INSTR_MEM[18]) );
  DFFR_X1 \INSTR_MEM_reg[17]  ( .D(n197), .CK(CLK), .RN(RST), .Q(INSTR_MEM[17]) );
  DFFR_X1 \INSTR_MEM_reg[16]  ( .D(n196), .CK(CLK), .RN(RST), .Q(INSTR_MEM[16]) );
  DFFR_X1 \INSTR_MEM_reg[15]  ( .D(n195), .CK(CLK), .RN(RST), .Q(INSTR_MEM[15]) );
  DFFR_X1 \INSTR_MEM_reg[14]  ( .D(n194), .CK(CLK), .RN(RST), .Q(INSTR_MEM[14]) );
  DFFR_X1 \INSTR_MEM_reg[13]  ( .D(n193), .CK(CLK), .RN(RST), .Q(INSTR_MEM[13]) );
  DFFR_X1 \INSTR_MEM_reg[12]  ( .D(n192), .CK(CLK), .RN(RST), .Q(INSTR_MEM[12]) );
  DFFR_X1 \INSTR_MEM_reg[11]  ( .D(n191), .CK(CLK), .RN(RST), .Q(INSTR_MEM[11]) );
  DFFR_X1 \CU_OUTS_WB_atMEM_reg[RF_WR_EN]  ( .D(n190), .CK(CLK), .RN(RST), .Q(
        \CU_OUTS_WB_atMEM[RF_WR_EN] ) );
  DFFR_X1 \CU_OUTS_MEM_atMEM_reg[DRAM_WR_EN][1]  ( .D(n189), .CK(CLK), .RN(RST), .Q(DRAM_WR_EN[1]) );
  DFFR_X1 \CU_OUTS_MEM_atMEM_reg[DRAM_WR_EN][0]  ( .D(n188), .CK(CLK), .RN(RST), .Q(DRAM_WR_EN[0]) );
  DFFR_X1 \INSTR_EXE_reg[31]  ( .D(n187), .CK(net18748), .RN(RST), .Q(
        INSTR_EXE[31]) );
  DFFR_X1 \INSTR_EXE_reg[29]  ( .D(n186), .CK(net18748), .RN(RST), .Q(
        INSTR_EXE[29]) );
  DFFR_X1 \INSTR_EXE_reg[27]  ( .D(n185), .CK(net18748), .RN(RST), .Q(
        INSTR_EXE[27]) );
  DFFR_X1 \INSTR_EXE_reg[20]  ( .D(n184), .CK(net18748), .RN(RST), .Q(
        INSTR_EXE[20]) );
  DFFR_X1 \INSTR_EXE_reg[19]  ( .D(n183), .CK(net18748), .RN(RST), .Q(
        INSTR_EXE[19]) );
  DFFR_X1 \INSTR_EXE_reg[18]  ( .D(n182), .CK(net18748), .RN(RST), .Q(
        INSTR_EXE[18]) );
  DFFR_X1 \INSTR_EXE_reg[17]  ( .D(n181), .CK(net18748), .RN(RST), .Q(
        INSTR_EXE[17]) );
  DFFR_X1 \INSTR_EXE_reg[16]  ( .D(n180), .CK(net18748), .RN(RST), .Q(
        INSTR_EXE[16]) );
  DFFR_X1 \INSTR_EXE_reg[15]  ( .D(n179), .CK(net18748), .RN(RST), .Q(
        INSTR_EXE[15]) );
  DFFR_X1 \INSTR_EXE_reg[14]  ( .D(n178), .CK(net18748), .RN(RST), .Q(
        INSTR_EXE[14]) );
  DFFR_X1 \INSTR_EXE_reg[13]  ( .D(n177), .CK(net18748), .RN(RST), .Q(
        INSTR_EXE[13]) );
  DFFR_X1 \INSTR_EXE_reg[12]  ( .D(n176), .CK(net18748), .RN(RST), .Q(
        INSTR_EXE[12]) );
  DFFR_X1 \INSTR_EXE_reg[11]  ( .D(n175), .CK(net18748), .RN(RST), .Q(
        INSTR_EXE[11]) );
  DFFR_X1 \INSTR_EXE_reg[5]  ( .D(n174), .CK(net18748), .RN(RST), .Q(
        INSTR_EXE[5]) );
  DFFR_X1 \INSTR_EXE_reg[4]  ( .D(n173), .CK(net18748), .RN(RST), .Q(
        INSTR_EXE[4]) );
  DFFR_X1 \INSTR_EXE_reg[3]  ( .D(n172), .CK(net18748), .RN(RST), .Q(
        INSTR_EXE[3]) );
  DFFR_X1 \INSTR_EXE_reg[2]  ( .D(n171), .CK(net18753), .RN(RST), .Q(
        INSTR_EXE[2]) );
  DFFR_X1 \INSTR_EXE_reg[1]  ( .D(n170), .CK(net18753), .RN(RST), .Q(
        INSTR_EXE[1]) );
  DFFR_X1 \INSTR_EXE_reg[0]  ( .D(n169), .CK(net18753), .RN(RST), .Q(
        INSTR_EXE[0]) );
  DFFR_X1 \CU_OUTS_MEM_atEXE_reg[DRAM_WR_EN][1]  ( .D(n168), .CK(net18753), 
        .RN(RST), .Q(\CU_OUTS_MEM_atEXE[DRAM_WR_EN][1] ) );
  DFFR_X1 \CU_OUTS_MEM_atEXE_reg[DRAM_WR_EN][0]  ( .D(n167), .CK(net18753), 
        .RN(RST), .Q(\CU_OUTS_MEM_atEXE[DRAM_WR_EN][0] ) );
  DFFR_X1 \CU_OUTS_EXE_atEXE_reg[MULT_EN]  ( .D(n166), .CK(net18753), .RN(RST), 
        .Q(\CU_OUTS_EXE_atEXE[MULT_EN] ) );
  DFFR_X1 \CU_OUTS_WB_atEXE_reg[RF_WR_EN]  ( .D(n165), .CK(net18753), .RN(RST), 
        .Q(\CU_OUTS_WB_atEXE[RF_WR_EN] ) );
  DFFR_X1 \INSTR_ID_reg[31]  ( .D(n164), .CK(net18743), .RN(RST), .Q(
        INSTR_ID[31]) );
  DFFR_X1 \INSTR_ID_reg[29]  ( .D(n163), .CK(net18743), .RN(RST), .Q(
        INSTR_ID[29]) );
  DFFR_X1 \INSTR_ID_reg[27]  ( .D(n162), .CK(net18743), .RN(RST), .Q(
        INSTR_ID[27]) );
  DFFR_X1 \INSTR_ID_reg[25]  ( .D(n161), .CK(net18743), .RN(RST), .Q(
        INSTR_ID[25]) );
  DFFR_X1 \INSTR_ID_reg[24]  ( .D(n160), .CK(net18743), .RN(RST), .Q(
        INSTR_ID[24]) );
  DFFR_X1 \INSTR_ID_reg[23]  ( .D(n159), .CK(net18743), .RN(RST), .Q(
        INSTR_ID[23]) );
  DFFR_X1 \INSTR_ID_reg[22]  ( .D(n158), .CK(net18743), .RN(RST), .Q(
        INSTR_ID[22]) );
  DFFR_X1 \INSTR_ID_reg[21]  ( .D(n157), .CK(net18743), .RN(RST), .Q(
        INSTR_ID[21]) );
  DFFR_X1 \INSTR_ID_reg[20]  ( .D(n156), .CK(net18743), .RN(RST), .Q(
        INSTR_ID[20]) );
  DFFR_X1 \INSTR_ID_reg[19]  ( .D(n155), .CK(net18743), .RN(RST), .Q(
        INSTR_ID[19]) );
  DFFR_X1 \INSTR_ID_reg[18]  ( .D(n154), .CK(net18743), .RN(RST), .Q(
        INSTR_ID[18]) );
  DFFR_X1 \INSTR_ID_reg[17]  ( .D(n153), .CK(net18743), .RN(RST), .Q(
        INSTR_ID[17]) );
  DFFR_X1 \INSTR_ID_reg[16]  ( .D(n152), .CK(net18743), .RN(RST), .Q(
        INSTR_ID[16]) );
  DFFR_X1 \INSTR_ID_reg[15]  ( .D(n151), .CK(net18743), .RN(RST), .Q(
        INSTR_ID[15]) );
  DFFR_X1 \INSTR_ID_reg[14]  ( .D(n150), .CK(net18743), .RN(RST), .Q(
        INSTR_ID[14]) );
  DFFR_X1 \INSTR_ID_reg[13]  ( .D(n149), .CK(net18743), .RN(RST), .Q(
        INSTR_ID[13]) );
  DFFR_X1 \INSTR_ID_reg[12]  ( .D(n148), .CK(net18743), .RN(RST), .Q(
        INSTR_ID[12]) );
  DFFR_X1 \INSTR_ID_reg[11]  ( .D(n147), .CK(net18743), .RN(RST), .Q(
        INSTR_ID[11]) );
  DFFR_X1 \INSTR_ID_reg[5]  ( .D(n146), .CK(net18743), .RN(RST), .Q(
        INSTR_ID[5]) );
  DFFR_X1 \INSTR_ID_reg[4]  ( .D(n145), .CK(net18743), .RN(RST), .Q(
        INSTR_ID[4]) );
  DFFR_X1 \INSTR_ID_reg[3]  ( .D(n144), .CK(net18743), .RN(RST), .Q(
        INSTR_ID[3]) );
  DFFR_X1 \INSTR_ID_reg[2]  ( .D(n143), .CK(net18743), .RN(RST), .Q(
        INSTR_ID[2]) );
  DFFR_X1 \INSTR_ID_reg[1]  ( .D(n142), .CK(net18743), .RN(RST), .Q(
        INSTR_ID[1]) );
  DFFR_X1 \INSTR_ID_reg[0]  ( .D(n141), .CK(net18743), .RN(RST), .Q(
        INSTR_ID[0]) );
  DFFS_X1 \CU_OUTS_EXE_atEXE_reg[ALU_OP][4]  ( .D(n210), .CK(net18753), .SN(
        RST), .QN(\CU_OUTS_EXE_atEXE[ALU_OP][4] ) );
  AND2_X1 U152 ( .A1(IRAM_OUT[0]), .A2(n204), .ZN(n141) );
  AND2_X1 U153 ( .A1(IRAM_OUT[1]), .A2(n204), .ZN(n142) );
  AND2_X1 U154 ( .A1(IRAM_OUT[2]), .A2(n204), .ZN(n143) );
  AND2_X1 U155 ( .A1(IRAM_OUT[3]), .A2(n204), .ZN(n144) );
  AND2_X1 U156 ( .A1(IRAM_OUT[4]), .A2(n204), .ZN(n145) );
  AND2_X1 U157 ( .A1(IRAM_OUT[5]), .A2(n204), .ZN(n146) );
  AND2_X1 U158 ( .A1(IRAM_OUT[11]), .A2(n204), .ZN(n147) );
  AND2_X1 U159 ( .A1(IRAM_OUT[12]), .A2(n204), .ZN(n148) );
  AND2_X1 U160 ( .A1(IRAM_OUT[13]), .A2(n204), .ZN(n149) );
  AND2_X1 U161 ( .A1(IRAM_OUT[14]), .A2(n204), .ZN(n150) );
  AND2_X1 U162 ( .A1(IRAM_OUT[15]), .A2(n204), .ZN(n151) );
  AND2_X1 U163 ( .A1(IRAM_OUT[16]), .A2(n204), .ZN(n152) );
  AND2_X1 U164 ( .A1(IRAM_OUT[17]), .A2(n204), .ZN(n153) );
  AND2_X1 U165 ( .A1(IRAM_OUT[18]), .A2(n204), .ZN(n154) );
  AND2_X1 U166 ( .A1(IRAM_OUT[19]), .A2(n204), .ZN(n155) );
  AND2_X1 U167 ( .A1(IRAM_OUT[20]), .A2(n204), .ZN(n156) );
  AND2_X1 U168 ( .A1(IRAM_OUT[21]), .A2(n204), .ZN(n157) );
  AND2_X1 U169 ( .A1(IRAM_OUT[22]), .A2(n204), .ZN(n158) );
  AND2_X1 U170 ( .A1(IRAM_OUT[23]), .A2(n204), .ZN(n159) );
  AND2_X1 U171 ( .A1(IRAM_OUT[24]), .A2(n204), .ZN(n160) );
  AND2_X1 U172 ( .A1(IRAM_OUT[25]), .A2(n204), .ZN(n161) );
  AND2_X1 U173 ( .A1(IRAM_OUT[27]), .A2(n204), .ZN(n162) );
  AND2_X1 U174 ( .A1(IRAM_OUT[29]), .A2(n204), .ZN(n163) );
  AND2_X1 U175 ( .A1(IRAM_OUT[31]), .A2(n204), .ZN(n164) );
  AND2_X1 U176 ( .A1(\CU_OUTS[WB][RF_WR_EN] ), .A2(n139), .ZN(n165) );
  AND2_X1 U177 ( .A1(\CU_OUTS[EXE][MULT_EN] ), .A2(n139), .ZN(n166) );
  AND2_X1 U178 ( .A1(\CU_OUTS[MEM][DRAM_WR_EN][0] ), .A2(n139), .ZN(n167) );
  AND2_X1 U179 ( .A1(\CU_OUTS[MEM][DRAM_WR_EN][1] ), .A2(n139), .ZN(n168) );
  AND2_X1 U180 ( .A1(INSTR_ID[0]), .A2(n139), .ZN(n169) );
  AND2_X1 U181 ( .A1(INSTR_ID[1]), .A2(n139), .ZN(n170) );
  AND2_X1 U182 ( .A1(INSTR_ID[2]), .A2(n139), .ZN(n171) );
  AND2_X1 U183 ( .A1(INSTR_ID[3]), .A2(n139), .ZN(n172) );
  AND2_X1 U184 ( .A1(INSTR_ID[4]), .A2(n139), .ZN(n173) );
  AND2_X1 U185 ( .A1(INSTR_ID[5]), .A2(n139), .ZN(n174) );
  AND2_X1 U186 ( .A1(INSTR_ID[11]), .A2(n139), .ZN(n175) );
  AND2_X1 U187 ( .A1(INSTR_ID[12]), .A2(n139), .ZN(n176) );
  AND2_X1 U188 ( .A1(INSTR_ID[13]), .A2(n139), .ZN(n177) );
  AND2_X1 U189 ( .A1(INSTR_ID[14]), .A2(n139), .ZN(n178) );
  AND2_X1 U190 ( .A1(INSTR_ID[15]), .A2(n139), .ZN(n179) );
  AND2_X1 U191 ( .A1(INSTR_ID[16]), .A2(n139), .ZN(n180) );
  AND2_X1 U192 ( .A1(INSTR_ID[17]), .A2(n139), .ZN(n181) );
  AND2_X1 U193 ( .A1(INSTR_ID[18]), .A2(n139), .ZN(n182) );
  AND2_X1 U194 ( .A1(INSTR_ID[19]), .A2(n139), .ZN(n183) );
  AND2_X1 U195 ( .A1(INSTR_ID[20]), .A2(n139), .ZN(n184) );
  AND2_X1 U196 ( .A1(INSTR_ID[27]), .A2(n139), .ZN(n185) );
  AND2_X1 U197 ( .A1(INSTR_ID[29]), .A2(n139), .ZN(n186) );
  AND2_X1 U198 ( .A1(INSTR_ID[31]), .A2(n139), .ZN(n187) );
  AND2_X1 U199 ( .A1(\CU_OUTS_MEM_atEXE[DRAM_WR_EN][0] ), .A2(n138), .ZN(n188)
         );
  AND2_X1 U200 ( .A1(\CU_OUTS_MEM_atEXE[DRAM_WR_EN][1] ), .A2(n138), .ZN(n189)
         );
  AND2_X1 U201 ( .A1(\CU_OUTS_WB_atEXE[RF_WR_EN] ), .A2(n138), .ZN(n190) );
  AND2_X1 U202 ( .A1(INSTR_EXE[11]), .A2(n138), .ZN(n191) );
  AND2_X1 U203 ( .A1(INSTR_EXE[12]), .A2(n138), .ZN(n192) );
  AND2_X1 U204 ( .A1(INSTR_EXE[13]), .A2(n138), .ZN(n193) );
  AND2_X1 U205 ( .A1(INSTR_EXE[14]), .A2(n138), .ZN(n194) );
  AND2_X1 U206 ( .A1(INSTR_EXE[15]), .A2(n138), .ZN(n195) );
  AND2_X1 U207 ( .A1(INSTR_EXE[16]), .A2(n138), .ZN(n196) );
  AND2_X1 U208 ( .A1(INSTR_EXE[17]), .A2(n138), .ZN(n197) );
  AND2_X1 U209 ( .A1(INSTR_EXE[18]), .A2(n138), .ZN(n198) );
  AND2_X1 U210 ( .A1(INSTR_EXE[19]), .A2(n138), .ZN(n199) );
  AND2_X1 U211 ( .A1(INSTR_EXE[20]), .A2(n138), .ZN(n200) );
  AND2_X1 U212 ( .A1(INSTR_EXE[27]), .A2(n138), .ZN(n201) );
  AND2_X1 U213 ( .A1(INSTR_EXE[29]), .A2(n138), .ZN(n202) );
  AND2_X1 U214 ( .A1(INSTR_EXE[31]), .A2(n138), .ZN(n203) );
  BUF_X2 U215 ( .A(n140), .Z(n204) );
  INV_X1 U216 ( .A(\HDU_OUTS[EXE_BUBBLE] ), .ZN(n139) );
  BUF_X1 U217 ( .A(\HDU_OUTS[ID_BUBBLE] ), .Z(n205) );
  INV_X1 U218 ( .A(\HDU_OUTS[MEM_BUBBLE] ), .ZN(n138) );
  NAND2_X1 U219 ( .A1(\CU_OUTS[EXE][ALU_OP][2] ), .A2(n139), .ZN(n206) );
  NAND2_X1 U220 ( .A1(\CU_OUTS[EXE][ALU_OP][0] ), .A2(n139), .ZN(n207) );
  NAND2_X1 U221 ( .A1(\CU_OUTS[EXE][ALU_OP][1] ), .A2(n139), .ZN(n208) );
  NAND2_X1 U222 ( .A1(\CU_OUTS[EXE][ALU_OP][3] ), .A2(n139), .ZN(n209) );
  NAND2_X1 U223 ( .A1(\CU_OUTS[EXE][ALU_OP][4] ), .A2(n139), .ZN(n210) );
  INV_X1 U224 ( .A(n215), .ZN(IRAM_ADDR[4]) );
  INV_X1 U225 ( .A(n216), .ZN(IRAM_ADDR[3]) );
  OR2_X1 U228 ( .A1(\HDU_OUTS[MEM_BUBBLE] ), .A2(INSTR_EXE[26]), .ZN(N100) );
  OR2_X1 U229 ( .A1(\HDU_OUTS[MEM_BUBBLE] ), .A2(INSTR_EXE[28]), .ZN(N102) );
  OR2_X1 U230 ( .A1(\HDU_OUTS[MEM_BUBBLE] ), .A2(INSTR_EXE[30]), .ZN(N104) );
  OR2_X1 U231 ( .A1(n205), .A2(IRAM_OUT[26]), .ZN(N32) );
  OR2_X1 U232 ( .A1(n205), .A2(IRAM_OUT[28]), .ZN(N34) );
  OR2_X1 U233 ( .A1(n205), .A2(IRAM_OUT[30]), .ZN(N36) );
  OR2_X1 U234 ( .A1(\HDU_OUTS[EXE_BUBBLE] ), .A2(\HDU_OUTS[ID_EN] ), .ZN(N39)
         );
  OR2_X1 U235 ( .A1(n205), .A2(\HDU_OUTS[IF_EN] ), .ZN(N5) );
  OR2_X1 U236 ( .A1(\HDU_OUTS[EXE_BUBBLE] ), .A2(INSTR_ID[26]), .ZN(N66) );
  OR2_X1 U237 ( .A1(\HDU_OUTS[EXE_BUBBLE] ), .A2(INSTR_ID[28]), .ZN(N68) );
  OR2_X1 U238 ( .A1(\HDU_OUTS[EXE_BUBBLE] ), .A2(INSTR_ID[30]), .ZN(N70) );
  INV_X1 U239 ( .A(\HDU_OUTS[ID_BUBBLE] ), .ZN(n140) );
endmodule

