package DRAM_package is	
	
	type DRAM_WR_EN_type is (
		DRAM_WR_OFF,
		DRAM_WR_B,
		DRAM_WR_H,
		DRAM_WR_W
	);
	
end package DRAM_package;