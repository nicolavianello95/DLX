library ieee; 
use ieee.std_logic_1164.all; 
use ieee.std_logic_unsigned.all;
use work.my_package.all;			--for XOR operator between a std_logic and a std_logic_vector

-- Top level module of the Pentium 4 adder
ENTITY  ADDER_P4 IS
	GENERIC (N_BIT	: integer := 32);	--number of bits. Must be a number from 4 to 32 and a multiple of 4
    PORT   (A		: in  std_logic_vector(N_BIT - 1 downto 0);		-- input operand 1
			B		: in  std_logic_vector(N_BIT - 1 downto 0);		-- input operand 2
			add_sub	: in  std_logic;								-- carry-in
			Cout	: out std_logic;								-- carry-out
			SUM		: out std_logic_vector(N_BIT -1 downto 0));		-- ouput sum
END ENTITY ADDER_P4;		

architecture STRUCTURAL of ADDER_P4 is

	component SUMGENERATOR IS
		GENERIC(Nblocks			: positive := 8;	--number of carry select block
				bits_per_block	: positive := 4);	--number of bit per each block
													--the number of input bits is equal to Nblocks*bits_per_block
		PORT (	A				: in  std_logic_vector(bits_per_block*Nblocks - 1 downto 0);	--data input 1
				B         		: in  std_logic_vector(bits_per_block*Nblocks - 1 downto 0);	--data input 2
				CARRY_SELECT	: in  std_logic_vector(Nblocks-1 downto 0);						--carries from sparse tree
				SUM				: out std_logic_vector(bits_per_block*Nblocks - 1 downto 0));	--data output
	end component; 
  
	component CARRY_GENERATOR IS
		GENERIC (Nbit	: positive := 32);								--number of bits for the structure. Must be between 4 and 32 and a multiple of 4
		PORT   (	A		: in  std_logic_vector(Nbit - 1 downto 0);	--input operand 1
					B		: in  std_logic_vector(Nbit - 1 downto 0);	--input operand 2
					Cin	: in  std_logic;								--carry-in
					Cout	: out std_logic_vector(Nbit/4 downto 0));	--carry-out generated by the tree
	end component; 
  
	signal tmp_co	: std_logic_vector(N_BIT/4	downto 0); -- used to connect the carries lines between the two modules
	signal B_xor	: std_logic_vector(N_BIT - 1 downto 0); -- B is changed if a subtraction incoming. If it is a sum, it doesn't change
BEGIN

	CLA_SPARSE_TREE: CARRY_GENERATOR 
		GENERIC MAP (Nbit => N_BIT)
		PORT MAP  (A => A,	B => B_xor, Cin	=> add_sub, Cout => tmp_co);

	CSA: SUMGENERATOR
		GENERIC MAP(Nblocks=> N_BIT/4, bits_per_block => 4)
		PORT MAP(A => A, B => B_xor , CARRY_SELECT => tmp_co (N_BIT/4-1 downto 0), SUM => SUM);
		 
	-- the most significant bit of the carries signal is the carry-out of the complete adder
	Cout <= tmp_co(N_BIT/4);
	
	-- Every bits of B pass through a xor gates with the Cin. In this way, when a subtraction arrives, Cin is set to 1
	-- so it complements bit by bit the input B. If arrives a sum, nothing change and the input B is simply copied 
	
	B_xor <= B xor add_sub;

end STRUCTURAL;

